// soc_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                                  //                               clk.clk
		input  wire [31:0] dcc_data_0_external_connection_export,    //    dcc_data_0_external_connection.export
		input  wire [31:0] dcc_data_10_external_connection_export,   //   dcc_data_10_external_connection.export
		input  wire [31:0] dcc_data_11_external_connection_export,   //   dcc_data_11_external_connection.export
		input  wire [31:0] dcc_data_12_external_connection_export,   //   dcc_data_12_external_connection.export
		input  wire [31:0] dcc_data_13_external_connection_export,   //   dcc_data_13_external_connection.export
		input  wire [31:0] dcc_data_14_external_connection_export,   //   dcc_data_14_external_connection.export
		input  wire [31:0] dcc_data_15_external_connection_export,   //   dcc_data_15_external_connection.export
		input  wire [31:0] dcc_data_16_external_connection_export,   //   dcc_data_16_external_connection.export
		input  wire [31:0] dcc_data_17_external_connection_export,   //   dcc_data_17_external_connection.export
		input  wire [31:0] dcc_data_18_external_connection_export,   //   dcc_data_18_external_connection.export
		input  wire [31:0] dcc_data_19_external_connection_export,   //   dcc_data_19_external_connection.export
		input  wire [31:0] dcc_data_1_external_connection_export,    //    dcc_data_1_external_connection.export
		input  wire [31:0] dcc_data_20_external_connection_export,   //   dcc_data_20_external_connection.export
		input  wire [31:0] dcc_data_21_external_connection_export,   //   dcc_data_21_external_connection.export
		input  wire [31:0] dcc_data_22_external_connection_export,   //   dcc_data_22_external_connection.export
		input  wire [31:0] dcc_data_23_external_connection_export,   //   dcc_data_23_external_connection.export
		input  wire [31:0] dcc_data_24_external_connection_export,   //   dcc_data_24_external_connection.export
		input  wire [31:0] dcc_data_25_external_connection_export,   //   dcc_data_25_external_connection.export
		input  wire [31:0] dcc_data_26_external_connection_export,   //   dcc_data_26_external_connection.export
		input  wire [31:0] dcc_data_27_external_connection_export,   //   dcc_data_27_external_connection.export
		input  wire [31:0] dcc_data_28_external_connection_export,   //   dcc_data_28_external_connection.export
		input  wire [31:0] dcc_data_29_external_connection_export,   //   dcc_data_29_external_connection.export
		input  wire [31:0] dcc_data_2_external_connection_export,    //    dcc_data_2_external_connection.export
		input  wire [31:0] dcc_data_30_external_connection_export,   //   dcc_data_30_external_connection.export
		input  wire [31:0] dcc_data_31_external_connection_export,   //   dcc_data_31_external_connection.export
		input  wire [31:0] dcc_data_3_external_connection_export,    //    dcc_data_3_external_connection.export
		input  wire [31:0] dcc_data_4_external_connection_export,    //    dcc_data_4_external_connection.export
		input  wire [31:0] dcc_data_5_external_connection_export,    //    dcc_data_5_external_connection.export
		input  wire [31:0] dcc_data_6_external_connection_export,    //    dcc_data_6_external_connection.export
		input  wire [31:0] dcc_data_7_external_connection_export,    //    dcc_data_7_external_connection.export
		input  wire [31:0] dcc_data_8_external_connection_export,    //    dcc_data_8_external_connection.export
		input  wire [31:0] dcc_data_9_external_connection_export,    //    dcc_data_9_external_connection.export
		input  wire [25:0] dcc_time_out_external_connection_export,  //  dcc_time_out_external_connection.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,         //          hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,        //         hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_dma_req0_dma_req,               //                hps_0_f2h_dma_req0.dma_req
		input  wire        hps_0_f2h_dma_req0_dma_single,            //                                  .dma_single
		output wire        hps_0_f2h_dma_req0_dma_ack,               //                                  .dma_ack
		input  wire        hps_0_f2h_dma_req1_dma_req,               //                hps_0_f2h_dma_req1.dma_req
		input  wire        hps_0_f2h_dma_req1_dma_single,            //                                  .dma_single
		output wire        hps_0_f2h_dma_req1_dma_ack,               //                                  .dma_ack
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,     //           hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,         //          hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,                  //                   hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,    //                      hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,      //                                  .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,      //                                  .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,      //                                  .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,      //                                  .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,      //                                  .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,      //                                  .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,       //                                  .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,    //                                  .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,    //                                  .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,    //                                  .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,      //                                  .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,      //                                  .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,      //                                  .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,        //                                  .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,        //                                  .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,        //                                  .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,        //                                  .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,        //                                  .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,        //                                  .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,        //                                  .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,         //                                  .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,         //                                  .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,        //                                  .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,         //                                  .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,         //                                  .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,         //                                  .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,         //                                  .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,         //                                  .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,         //                                  .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,         //                                  .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,         //                                  .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,         //                                  .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,         //                                  .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,        //                                  .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,        //                                  .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,        //                                  .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,        //                                  .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim0_inst_CLK,       //                                  .hps_io_spim0_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim0_inst_MOSI,      //                                  .hps_io_spim0_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim0_inst_MISO,      //                                  .hps_io_spim0_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim0_inst_SS0,       //                                  .hps_io_spim0_inst_SS0
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,       //                                  .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,      //                                  .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,      //                                  .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,       //                                  .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,        //                                  .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,        //                                  .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,        //                                  .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,        //                                  .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,        //                                  .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,        //                                  .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,     //                                  .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,     //                                  .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO37,     //                                  .hps_io_gpio_inst_GPIO37
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,     //                                  .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,     //                                  .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO44,     //                                  .hps_io_gpio_inst_GPIO44
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,     //                                  .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,     //                                  .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,     //                                  .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,     //                                  .hps_io_gpio_inst_GPIO61
		output wire        hps_read_bit_external_connection_export,  //  hps_read_bit_external_connection.export
		output wire [9:0]  ledr_external_connection_export,          //          ledr_external_connection.export
		output wire [14:0] memory_mem_a,                             //                            memory.mem_a
		output wire [2:0]  memory_mem_ba,                            //                                  .mem_ba
		output wire        memory_mem_ck,                            //                                  .mem_ck
		output wire        memory_mem_ck_n,                          //                                  .mem_ck_n
		output wire        memory_mem_cke,                           //                                  .mem_cke
		output wire        memory_mem_cs_n,                          //                                  .mem_cs_n
		output wire        memory_mem_ras_n,                         //                                  .mem_ras_n
		output wire        memory_mem_cas_n,                         //                                  .mem_cas_n
		output wire        memory_mem_we_n,                          //                                  .mem_we_n
		output wire        memory_mem_reset_n,                       //                                  .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                            //                                  .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                           //                                  .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                         //                                  .mem_dqs_n
		output wire        memory_mem_odt,                           //                                  .mem_odt
		output wire [3:0]  memory_mem_dm,                            //                                  .mem_dm
		input  wire        memory_oct_rzqin,                         //                                  .oct_rzqin
		input  wire [31:0] pps_count_out_external_connection_export, // pps_count_out_external_connection.export
		input  wire        reset_reset_n,                            //                             reset.reset_n
		input  wire [13:0] sw_external_connection_export             //            sw_external_connection.export
	);

	wire  [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [17:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire         mm_bridge_0_m0_waitrequest;                                // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [31:0] mm_bridge_0_m0_readdata;                                   // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire  [17:0] mm_bridge_0_m0_address;                                    // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire         mm_bridge_0_m0_read;                                       // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire   [3:0] mm_bridge_0_m0_byteenable;                                 // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                              // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire  [31:0] mm_bridge_0_m0_writedata;                                  // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                      // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire   [0:0] mm_bridge_0_m0_burstcount;                                 // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire  [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [17:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [63:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [7:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [63:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                      // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                        // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                         // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                           // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                       // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_0_sw_s1_chipselect;                        // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                           // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_sw_s1_write;                             // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                         // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_0_dcc_data_0_s1_chipselect;                // mm_interconnect_0:dcc_data_0_s1_chipselect -> dcc_data_0:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_0_s1_readdata;                  // dcc_data_0:readdata -> mm_interconnect_0:dcc_data_0_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_0_s1_address;                   // mm_interconnect_0:dcc_data_0_s1_address -> dcc_data_0:address
	wire         mm_interconnect_0_dcc_data_0_s1_write;                     // mm_interconnect_0:dcc_data_0_s1_write -> dcc_data_0:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_0_s1_writedata;                 // mm_interconnect_0:dcc_data_0_s1_writedata -> dcc_data_0:writedata
	wire         mm_interconnect_0_hps_read_bit_s1_chipselect;              // mm_interconnect_0:hps_read_bit_s1_chipselect -> hps_read_bit:chipselect
	wire  [31:0] mm_interconnect_0_hps_read_bit_s1_readdata;                // hps_read_bit:readdata -> mm_interconnect_0:hps_read_bit_s1_readdata
	wire   [1:0] mm_interconnect_0_hps_read_bit_s1_address;                 // mm_interconnect_0:hps_read_bit_s1_address -> hps_read_bit:address
	wire         mm_interconnect_0_hps_read_bit_s1_write;                   // mm_interconnect_0:hps_read_bit_s1_write -> hps_read_bit:write_n
	wire  [31:0] mm_interconnect_0_hps_read_bit_s1_writedata;               // mm_interconnect_0:hps_read_bit_s1_writedata -> hps_read_bit:writedata
	wire         mm_interconnect_0_dcc_data_1_s1_chipselect;                // mm_interconnect_0:dcc_data_1_s1_chipselect -> dcc_data_1:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_1_s1_readdata;                  // dcc_data_1:readdata -> mm_interconnect_0:dcc_data_1_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_1_s1_address;                   // mm_interconnect_0:dcc_data_1_s1_address -> dcc_data_1:address
	wire         mm_interconnect_0_dcc_data_1_s1_write;                     // mm_interconnect_0:dcc_data_1_s1_write -> dcc_data_1:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_1_s1_writedata;                 // mm_interconnect_0:dcc_data_1_s1_writedata -> dcc_data_1:writedata
	wire         mm_interconnect_0_dcc_time_out_s1_chipselect;              // mm_interconnect_0:dcc_time_out_s1_chipselect -> dcc_time_out:chipselect
	wire  [31:0] mm_interconnect_0_dcc_time_out_s1_readdata;                // dcc_time_out:readdata -> mm_interconnect_0:dcc_time_out_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_time_out_s1_address;                 // mm_interconnect_0:dcc_time_out_s1_address -> dcc_time_out:address
	wire         mm_interconnect_0_dcc_time_out_s1_write;                   // mm_interconnect_0:dcc_time_out_s1_write -> dcc_time_out:write_n
	wire  [31:0] mm_interconnect_0_dcc_time_out_s1_writedata;               // mm_interconnect_0:dcc_time_out_s1_writedata -> dcc_time_out:writedata
	wire         mm_interconnect_0_dcc_data_2_s1_chipselect;                // mm_interconnect_0:dcc_data_2_s1_chipselect -> dcc_data_2:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_2_s1_readdata;                  // dcc_data_2:readdata -> mm_interconnect_0:dcc_data_2_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_2_s1_address;                   // mm_interconnect_0:dcc_data_2_s1_address -> dcc_data_2:address
	wire         mm_interconnect_0_dcc_data_2_s1_write;                     // mm_interconnect_0:dcc_data_2_s1_write -> dcc_data_2:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_2_s1_writedata;                 // mm_interconnect_0:dcc_data_2_s1_writedata -> dcc_data_2:writedata
	wire         mm_interconnect_0_dcc_data_3_s1_chipselect;                // mm_interconnect_0:dcc_data_3_s1_chipselect -> dcc_data_3:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_3_s1_readdata;                  // dcc_data_3:readdata -> mm_interconnect_0:dcc_data_3_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_3_s1_address;                   // mm_interconnect_0:dcc_data_3_s1_address -> dcc_data_3:address
	wire         mm_interconnect_0_dcc_data_3_s1_write;                     // mm_interconnect_0:dcc_data_3_s1_write -> dcc_data_3:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_3_s1_writedata;                 // mm_interconnect_0:dcc_data_3_s1_writedata -> dcc_data_3:writedata
	wire         mm_interconnect_0_dcc_data_4_s1_chipselect;                // mm_interconnect_0:dcc_data_4_s1_chipselect -> dcc_data_4:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_4_s1_readdata;                  // dcc_data_4:readdata -> mm_interconnect_0:dcc_data_4_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_4_s1_address;                   // mm_interconnect_0:dcc_data_4_s1_address -> dcc_data_4:address
	wire         mm_interconnect_0_dcc_data_4_s1_write;                     // mm_interconnect_0:dcc_data_4_s1_write -> dcc_data_4:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_4_s1_writedata;                 // mm_interconnect_0:dcc_data_4_s1_writedata -> dcc_data_4:writedata
	wire         mm_interconnect_0_dcc_data_5_s1_chipselect;                // mm_interconnect_0:dcc_data_5_s1_chipselect -> dcc_data_5:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_5_s1_readdata;                  // dcc_data_5:readdata -> mm_interconnect_0:dcc_data_5_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_5_s1_address;                   // mm_interconnect_0:dcc_data_5_s1_address -> dcc_data_5:address
	wire         mm_interconnect_0_dcc_data_5_s1_write;                     // mm_interconnect_0:dcc_data_5_s1_write -> dcc_data_5:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_5_s1_writedata;                 // mm_interconnect_0:dcc_data_5_s1_writedata -> dcc_data_5:writedata
	wire         mm_interconnect_0_dcc_data_6_s1_chipselect;                // mm_interconnect_0:dcc_data_6_s1_chipselect -> dcc_data_6:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_6_s1_readdata;                  // dcc_data_6:readdata -> mm_interconnect_0:dcc_data_6_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_6_s1_address;                   // mm_interconnect_0:dcc_data_6_s1_address -> dcc_data_6:address
	wire         mm_interconnect_0_dcc_data_6_s1_write;                     // mm_interconnect_0:dcc_data_6_s1_write -> dcc_data_6:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_6_s1_writedata;                 // mm_interconnect_0:dcc_data_6_s1_writedata -> dcc_data_6:writedata
	wire         mm_interconnect_0_dcc_data_7_s1_chipselect;                // mm_interconnect_0:dcc_data_7_s1_chipselect -> dcc_data_7:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_7_s1_readdata;                  // dcc_data_7:readdata -> mm_interconnect_0:dcc_data_7_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_7_s1_address;                   // mm_interconnect_0:dcc_data_7_s1_address -> dcc_data_7:address
	wire         mm_interconnect_0_dcc_data_7_s1_write;                     // mm_interconnect_0:dcc_data_7_s1_write -> dcc_data_7:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_7_s1_writedata;                 // mm_interconnect_0:dcc_data_7_s1_writedata -> dcc_data_7:writedata
	wire         mm_interconnect_0_dcc_data_8_s1_chipselect;                // mm_interconnect_0:dcc_data_8_s1_chipselect -> dcc_data_8:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_8_s1_readdata;                  // dcc_data_8:readdata -> mm_interconnect_0:dcc_data_8_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_8_s1_address;                   // mm_interconnect_0:dcc_data_8_s1_address -> dcc_data_8:address
	wire         mm_interconnect_0_dcc_data_8_s1_write;                     // mm_interconnect_0:dcc_data_8_s1_write -> dcc_data_8:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_8_s1_writedata;                 // mm_interconnect_0:dcc_data_8_s1_writedata -> dcc_data_8:writedata
	wire         mm_interconnect_0_dcc_data_9_s1_chipselect;                // mm_interconnect_0:dcc_data_9_s1_chipselect -> dcc_data_9:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_9_s1_readdata;                  // dcc_data_9:readdata -> mm_interconnect_0:dcc_data_9_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_9_s1_address;                   // mm_interconnect_0:dcc_data_9_s1_address -> dcc_data_9:address
	wire         mm_interconnect_0_dcc_data_9_s1_write;                     // mm_interconnect_0:dcc_data_9_s1_write -> dcc_data_9:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_9_s1_writedata;                 // mm_interconnect_0:dcc_data_9_s1_writedata -> dcc_data_9:writedata
	wire         mm_interconnect_0_dcc_data_10_s1_chipselect;               // mm_interconnect_0:dcc_data_10_s1_chipselect -> dcc_data_10:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_10_s1_readdata;                 // dcc_data_10:readdata -> mm_interconnect_0:dcc_data_10_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_10_s1_address;                  // mm_interconnect_0:dcc_data_10_s1_address -> dcc_data_10:address
	wire         mm_interconnect_0_dcc_data_10_s1_write;                    // mm_interconnect_0:dcc_data_10_s1_write -> dcc_data_10:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_10_s1_writedata;                // mm_interconnect_0:dcc_data_10_s1_writedata -> dcc_data_10:writedata
	wire         mm_interconnect_0_dcc_data_11_s1_chipselect;               // mm_interconnect_0:dcc_data_11_s1_chipselect -> dcc_data_11:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_11_s1_readdata;                 // dcc_data_11:readdata -> mm_interconnect_0:dcc_data_11_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_11_s1_address;                  // mm_interconnect_0:dcc_data_11_s1_address -> dcc_data_11:address
	wire         mm_interconnect_0_dcc_data_11_s1_write;                    // mm_interconnect_0:dcc_data_11_s1_write -> dcc_data_11:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_11_s1_writedata;                // mm_interconnect_0:dcc_data_11_s1_writedata -> dcc_data_11:writedata
	wire         mm_interconnect_0_dcc_data_12_s1_chipselect;               // mm_interconnect_0:dcc_data_12_s1_chipselect -> dcc_data_12:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_12_s1_readdata;                 // dcc_data_12:readdata -> mm_interconnect_0:dcc_data_12_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_12_s1_address;                  // mm_interconnect_0:dcc_data_12_s1_address -> dcc_data_12:address
	wire         mm_interconnect_0_dcc_data_12_s1_write;                    // mm_interconnect_0:dcc_data_12_s1_write -> dcc_data_12:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_12_s1_writedata;                // mm_interconnect_0:dcc_data_12_s1_writedata -> dcc_data_12:writedata
	wire         mm_interconnect_0_dcc_data_13_s1_chipselect;               // mm_interconnect_0:dcc_data_13_s1_chipselect -> dcc_data_13:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_13_s1_readdata;                 // dcc_data_13:readdata -> mm_interconnect_0:dcc_data_13_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_13_s1_address;                  // mm_interconnect_0:dcc_data_13_s1_address -> dcc_data_13:address
	wire         mm_interconnect_0_dcc_data_13_s1_write;                    // mm_interconnect_0:dcc_data_13_s1_write -> dcc_data_13:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_13_s1_writedata;                // mm_interconnect_0:dcc_data_13_s1_writedata -> dcc_data_13:writedata
	wire         mm_interconnect_0_dcc_data_14_s1_chipselect;               // mm_interconnect_0:dcc_data_14_s1_chipselect -> dcc_data_14:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_14_s1_readdata;                 // dcc_data_14:readdata -> mm_interconnect_0:dcc_data_14_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_14_s1_address;                  // mm_interconnect_0:dcc_data_14_s1_address -> dcc_data_14:address
	wire         mm_interconnect_0_dcc_data_14_s1_write;                    // mm_interconnect_0:dcc_data_14_s1_write -> dcc_data_14:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_14_s1_writedata;                // mm_interconnect_0:dcc_data_14_s1_writedata -> dcc_data_14:writedata
	wire         mm_interconnect_0_dcc_data_15_s1_chipselect;               // mm_interconnect_0:dcc_data_15_s1_chipselect -> dcc_data_15:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_15_s1_readdata;                 // dcc_data_15:readdata -> mm_interconnect_0:dcc_data_15_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_15_s1_address;                  // mm_interconnect_0:dcc_data_15_s1_address -> dcc_data_15:address
	wire         mm_interconnect_0_dcc_data_15_s1_write;                    // mm_interconnect_0:dcc_data_15_s1_write -> dcc_data_15:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_15_s1_writedata;                // mm_interconnect_0:dcc_data_15_s1_writedata -> dcc_data_15:writedata
	wire         mm_interconnect_0_dcc_data_16_s1_chipselect;               // mm_interconnect_0:dcc_data_16_s1_chipselect -> dcc_data_16:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_16_s1_readdata;                 // dcc_data_16:readdata -> mm_interconnect_0:dcc_data_16_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_16_s1_address;                  // mm_interconnect_0:dcc_data_16_s1_address -> dcc_data_16:address
	wire         mm_interconnect_0_dcc_data_16_s1_write;                    // mm_interconnect_0:dcc_data_16_s1_write -> dcc_data_16:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_16_s1_writedata;                // mm_interconnect_0:dcc_data_16_s1_writedata -> dcc_data_16:writedata
	wire         mm_interconnect_0_dcc_data_17_s1_chipselect;               // mm_interconnect_0:dcc_data_17_s1_chipselect -> dcc_data_17:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_17_s1_readdata;                 // dcc_data_17:readdata -> mm_interconnect_0:dcc_data_17_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_17_s1_address;                  // mm_interconnect_0:dcc_data_17_s1_address -> dcc_data_17:address
	wire         mm_interconnect_0_dcc_data_17_s1_write;                    // mm_interconnect_0:dcc_data_17_s1_write -> dcc_data_17:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_17_s1_writedata;                // mm_interconnect_0:dcc_data_17_s1_writedata -> dcc_data_17:writedata
	wire         mm_interconnect_0_dcc_data_18_s1_chipselect;               // mm_interconnect_0:dcc_data_18_s1_chipselect -> dcc_data_18:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_18_s1_readdata;                 // dcc_data_18:readdata -> mm_interconnect_0:dcc_data_18_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_18_s1_address;                  // mm_interconnect_0:dcc_data_18_s1_address -> dcc_data_18:address
	wire         mm_interconnect_0_dcc_data_18_s1_write;                    // mm_interconnect_0:dcc_data_18_s1_write -> dcc_data_18:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_18_s1_writedata;                // mm_interconnect_0:dcc_data_18_s1_writedata -> dcc_data_18:writedata
	wire         mm_interconnect_0_dcc_data_19_s1_chipselect;               // mm_interconnect_0:dcc_data_19_s1_chipselect -> dcc_data_19:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_19_s1_readdata;                 // dcc_data_19:readdata -> mm_interconnect_0:dcc_data_19_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_19_s1_address;                  // mm_interconnect_0:dcc_data_19_s1_address -> dcc_data_19:address
	wire         mm_interconnect_0_dcc_data_19_s1_write;                    // mm_interconnect_0:dcc_data_19_s1_write -> dcc_data_19:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_19_s1_writedata;                // mm_interconnect_0:dcc_data_19_s1_writedata -> dcc_data_19:writedata
	wire         mm_interconnect_0_dcc_data_20_s1_chipselect;               // mm_interconnect_0:dcc_data_20_s1_chipselect -> dcc_data_20:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_20_s1_readdata;                 // dcc_data_20:readdata -> mm_interconnect_0:dcc_data_20_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_20_s1_address;                  // mm_interconnect_0:dcc_data_20_s1_address -> dcc_data_20:address
	wire         mm_interconnect_0_dcc_data_20_s1_write;                    // mm_interconnect_0:dcc_data_20_s1_write -> dcc_data_20:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_20_s1_writedata;                // mm_interconnect_0:dcc_data_20_s1_writedata -> dcc_data_20:writedata
	wire         mm_interconnect_0_dcc_data_21_s1_chipselect;               // mm_interconnect_0:dcc_data_21_s1_chipselect -> dcc_data_21:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_21_s1_readdata;                 // dcc_data_21:readdata -> mm_interconnect_0:dcc_data_21_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_21_s1_address;                  // mm_interconnect_0:dcc_data_21_s1_address -> dcc_data_21:address
	wire         mm_interconnect_0_dcc_data_21_s1_write;                    // mm_interconnect_0:dcc_data_21_s1_write -> dcc_data_21:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_21_s1_writedata;                // mm_interconnect_0:dcc_data_21_s1_writedata -> dcc_data_21:writedata
	wire         mm_interconnect_0_dcc_data_22_s1_chipselect;               // mm_interconnect_0:dcc_data_22_s1_chipselect -> dcc_data_22:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_22_s1_readdata;                 // dcc_data_22:readdata -> mm_interconnect_0:dcc_data_22_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_22_s1_address;                  // mm_interconnect_0:dcc_data_22_s1_address -> dcc_data_22:address
	wire         mm_interconnect_0_dcc_data_22_s1_write;                    // mm_interconnect_0:dcc_data_22_s1_write -> dcc_data_22:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_22_s1_writedata;                // mm_interconnect_0:dcc_data_22_s1_writedata -> dcc_data_22:writedata
	wire         mm_interconnect_0_dcc_data_23_s1_chipselect;               // mm_interconnect_0:dcc_data_23_s1_chipselect -> dcc_data_23:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_23_s1_readdata;                 // dcc_data_23:readdata -> mm_interconnect_0:dcc_data_23_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_23_s1_address;                  // mm_interconnect_0:dcc_data_23_s1_address -> dcc_data_23:address
	wire         mm_interconnect_0_dcc_data_23_s1_write;                    // mm_interconnect_0:dcc_data_23_s1_write -> dcc_data_23:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_23_s1_writedata;                // mm_interconnect_0:dcc_data_23_s1_writedata -> dcc_data_23:writedata
	wire         mm_interconnect_0_dcc_data_24_s1_chipselect;               // mm_interconnect_0:dcc_data_24_s1_chipselect -> dcc_data_24:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_24_s1_readdata;                 // dcc_data_24:readdata -> mm_interconnect_0:dcc_data_24_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_24_s1_address;                  // mm_interconnect_0:dcc_data_24_s1_address -> dcc_data_24:address
	wire         mm_interconnect_0_dcc_data_24_s1_write;                    // mm_interconnect_0:dcc_data_24_s1_write -> dcc_data_24:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_24_s1_writedata;                // mm_interconnect_0:dcc_data_24_s1_writedata -> dcc_data_24:writedata
	wire         mm_interconnect_0_dcc_data_25_s1_chipselect;               // mm_interconnect_0:dcc_data_25_s1_chipselect -> dcc_data_25:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_25_s1_readdata;                 // dcc_data_25:readdata -> mm_interconnect_0:dcc_data_25_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_25_s1_address;                  // mm_interconnect_0:dcc_data_25_s1_address -> dcc_data_25:address
	wire         mm_interconnect_0_dcc_data_25_s1_write;                    // mm_interconnect_0:dcc_data_25_s1_write -> dcc_data_25:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_25_s1_writedata;                // mm_interconnect_0:dcc_data_25_s1_writedata -> dcc_data_25:writedata
	wire         mm_interconnect_0_dcc_data_26_s1_chipselect;               // mm_interconnect_0:dcc_data_26_s1_chipselect -> dcc_data_26:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_26_s1_readdata;                 // dcc_data_26:readdata -> mm_interconnect_0:dcc_data_26_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_26_s1_address;                  // mm_interconnect_0:dcc_data_26_s1_address -> dcc_data_26:address
	wire         mm_interconnect_0_dcc_data_26_s1_write;                    // mm_interconnect_0:dcc_data_26_s1_write -> dcc_data_26:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_26_s1_writedata;                // mm_interconnect_0:dcc_data_26_s1_writedata -> dcc_data_26:writedata
	wire         mm_interconnect_0_dcc_data_27_s1_chipselect;               // mm_interconnect_0:dcc_data_27_s1_chipselect -> dcc_data_27:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_27_s1_readdata;                 // dcc_data_27:readdata -> mm_interconnect_0:dcc_data_27_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_27_s1_address;                  // mm_interconnect_0:dcc_data_27_s1_address -> dcc_data_27:address
	wire         mm_interconnect_0_dcc_data_27_s1_write;                    // mm_interconnect_0:dcc_data_27_s1_write -> dcc_data_27:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_27_s1_writedata;                // mm_interconnect_0:dcc_data_27_s1_writedata -> dcc_data_27:writedata
	wire         mm_interconnect_0_dcc_data_28_s1_chipselect;               // mm_interconnect_0:dcc_data_28_s1_chipselect -> dcc_data_28:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_28_s1_readdata;                 // dcc_data_28:readdata -> mm_interconnect_0:dcc_data_28_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_28_s1_address;                  // mm_interconnect_0:dcc_data_28_s1_address -> dcc_data_28:address
	wire         mm_interconnect_0_dcc_data_28_s1_write;                    // mm_interconnect_0:dcc_data_28_s1_write -> dcc_data_28:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_28_s1_writedata;                // mm_interconnect_0:dcc_data_28_s1_writedata -> dcc_data_28:writedata
	wire         mm_interconnect_0_dcc_data_29_s1_chipselect;               // mm_interconnect_0:dcc_data_29_s1_chipselect -> dcc_data_29:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_29_s1_readdata;                 // dcc_data_29:readdata -> mm_interconnect_0:dcc_data_29_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_29_s1_address;                  // mm_interconnect_0:dcc_data_29_s1_address -> dcc_data_29:address
	wire         mm_interconnect_0_dcc_data_29_s1_write;                    // mm_interconnect_0:dcc_data_29_s1_write -> dcc_data_29:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_29_s1_writedata;                // mm_interconnect_0:dcc_data_29_s1_writedata -> dcc_data_29:writedata
	wire         mm_interconnect_0_dcc_data_30_s1_chipselect;               // mm_interconnect_0:dcc_data_30_s1_chipselect -> dcc_data_30:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_30_s1_readdata;                 // dcc_data_30:readdata -> mm_interconnect_0:dcc_data_30_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_30_s1_address;                  // mm_interconnect_0:dcc_data_30_s1_address -> dcc_data_30:address
	wire         mm_interconnect_0_dcc_data_30_s1_write;                    // mm_interconnect_0:dcc_data_30_s1_write -> dcc_data_30:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_30_s1_writedata;                // mm_interconnect_0:dcc_data_30_s1_writedata -> dcc_data_30:writedata
	wire         mm_interconnect_0_dcc_data_31_s1_chipselect;               // mm_interconnect_0:dcc_data_31_s1_chipselect -> dcc_data_31:chipselect
	wire  [31:0] mm_interconnect_0_dcc_data_31_s1_readdata;                 // dcc_data_31:readdata -> mm_interconnect_0:dcc_data_31_s1_readdata
	wire   [1:0] mm_interconnect_0_dcc_data_31_s1_address;                  // mm_interconnect_0:dcc_data_31_s1_address -> dcc_data_31:address
	wire         mm_interconnect_0_dcc_data_31_s1_write;                    // mm_interconnect_0:dcc_data_31_s1_write -> dcc_data_31:write_n
	wire  [31:0] mm_interconnect_0_dcc_data_31_s1_writedata;                // mm_interconnect_0:dcc_data_31_s1_writedata -> dcc_data_31:writedata
	wire         mm_interconnect_0_pps_count_out_s1_chipselect;             // mm_interconnect_0:pps_count_out_s1_chipselect -> pps_count_out:chipselect
	wire  [31:0] mm_interconnect_0_pps_count_out_s1_readdata;               // pps_count_out:readdata -> mm_interconnect_0:pps_count_out_s1_readdata
	wire   [1:0] mm_interconnect_0_pps_count_out_s1_address;                // mm_interconnect_0:pps_count_out_s1_address -> pps_count_out:address
	wire         mm_interconnect_0_pps_count_out_s1_write;                  // mm_interconnect_0:pps_count_out_s1_write -> pps_count_out:write_n
	wire  [31:0] mm_interconnect_0_pps_count_out_s1_writedata;              // mm_interconnect_0:pps_count_out_s1_writedata -> pps_count_out:writedata
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                           // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                             // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                             // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                            // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                             // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                               // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                           // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                            // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                            // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                            // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                            // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                             // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                           // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                           // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                              // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                            // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                            // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                            // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                           // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                            // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                            // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                             // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                             // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                              // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                            // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                           // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                            // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_readdata;                 // mm_bridge_0:s0_readdata -> mm_interconnect_1:mm_bridge_0_s0_readdata
	wire         mm_interconnect_1_mm_bridge_0_s0_waitrequest;              // mm_bridge_0:s0_waitrequest -> mm_interconnect_1:mm_bridge_0_s0_waitrequest
	wire         mm_interconnect_1_mm_bridge_0_s0_debugaccess;              // mm_interconnect_1:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire  [17:0] mm_interconnect_1_mm_bridge_0_s0_address;                  // mm_interconnect_1:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_1_mm_bridge_0_s0_read;                     // mm_interconnect_1:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire   [3:0] mm_interconnect_1_mm_bridge_0_s0_byteenable;               // mm_interconnect_1:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_1_mm_bridge_0_s0_readdatavalid;            // mm_bridge_0:s0_readdatavalid -> mm_interconnect_1:mm_bridge_0_s0_readdatavalid
	wire         mm_interconnect_1_mm_bridge_0_s0_write;                    // mm_interconnect_1:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_writedata;                // mm_interconnect_1:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_1_mm_bridge_0_s0_burstcount;               // mm_interconnect_1:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire         irq_mapper_receiver0_irq;                                  // sw:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // dcc_data_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // dcc_data_1:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // dcc_time_out:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // dcc_data_2:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // dcc_data_3:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                  // dcc_data_4:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                  // dcc_data_5:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                  // dcc_data_6:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                  // dcc_data_7:irq -> irq_mapper:receiver9_irq
	wire         irq_mapper_receiver10_irq;                                 // dcc_data_8:irq -> irq_mapper:receiver10_irq
	wire         irq_mapper_receiver11_irq;                                 // dcc_data_9:irq -> irq_mapper:receiver11_irq
	wire         irq_mapper_receiver12_irq;                                 // dcc_data_10:irq -> irq_mapper:receiver12_irq
	wire         irq_mapper_receiver13_irq;                                 // dcc_data_11:irq -> irq_mapper:receiver13_irq
	wire         irq_mapper_receiver14_irq;                                 // dcc_data_12:irq -> irq_mapper:receiver14_irq
	wire         irq_mapper_receiver15_irq;                                 // dcc_data_13:irq -> irq_mapper:receiver15_irq
	wire         irq_mapper_receiver16_irq;                                 // dcc_data_14:irq -> irq_mapper:receiver16_irq
	wire         irq_mapper_receiver17_irq;                                 // dcc_data_15:irq -> irq_mapper:receiver17_irq
	wire         irq_mapper_receiver18_irq;                                 // pps_count_out:irq -> irq_mapper:receiver18_irq
	wire  [31:0] hps_0_f2h_irq0_irq;                                        // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire         irq_mapper_001_receiver0_irq;                              // dcc_data_17:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                              // dcc_data_18:irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver2_irq;                              // dcc_data_19:irq -> irq_mapper_001:receiver2_irq
	wire         irq_mapper_001_receiver3_irq;                              // dcc_data_20:irq -> irq_mapper_001:receiver3_irq
	wire         irq_mapper_001_receiver4_irq;                              // dcc_data_21:irq -> irq_mapper_001:receiver4_irq
	wire         irq_mapper_001_receiver5_irq;                              // dcc_data_22:irq -> irq_mapper_001:receiver5_irq
	wire         irq_mapper_001_receiver6_irq;                              // dcc_data_23:irq -> irq_mapper_001:receiver6_irq
	wire         irq_mapper_001_receiver7_irq;                              // dcc_data_24:irq -> irq_mapper_001:receiver7_irq
	wire         irq_mapper_001_receiver8_irq;                              // dcc_data_25:irq -> irq_mapper_001:receiver8_irq
	wire         irq_mapper_001_receiver9_irq;                              // dcc_data_26:irq -> irq_mapper_001:receiver9_irq
	wire         irq_mapper_001_receiver10_irq;                             // dcc_data_27:irq -> irq_mapper_001:receiver10_irq
	wire         irq_mapper_001_receiver11_irq;                             // dcc_data_28:irq -> irq_mapper_001:receiver11_irq
	wire         irq_mapper_001_receiver12_irq;                             // dcc_data_29:irq -> irq_mapper_001:receiver12_irq
	wire         irq_mapper_001_receiver13_irq;                             // dcc_data_30:irq -> irq_mapper_001:receiver13_irq
	wire         irq_mapper_001_receiver14_irq;                             // dcc_data_31:irq -> irq_mapper_001:receiver14_irq
	wire         irq_mapper_001_receiver15_irq;                             // dcc_data_16:irq -> irq_mapper_001:receiver15_irq
	wire  [31:0] hps_0_f2h_irq1_irq;                                        // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         irq_mapper_002_receiver0_irq;                              // timer:irq -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                              // jtag_uart:av_irq -> irq_mapper_002:receiver1_irq
	wire  [31:0] nios2_gen2_irq_irq;                                        // irq_mapper_002:sender_irq -> nios2_gen2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [dcc_data_0:reset_n, dcc_data_10:reset_n, dcc_data_11:reset_n, dcc_data_12:reset_n, dcc_data_13:reset_n, dcc_data_14:reset_n, dcc_data_15:reset_n, dcc_data_16:reset_n, dcc_data_17:reset_n, dcc_data_18:reset_n, dcc_data_19:reset_n, dcc_data_1:reset_n, dcc_data_20:reset_n, dcc_data_21:reset_n, dcc_data_22:reset_n, dcc_data_23:reset_n, dcc_data_24:reset_n, dcc_data_25:reset_n, dcc_data_26:reset_n, dcc_data_27:reset_n, dcc_data_28:reset_n, dcc_data_29:reset_n, dcc_data_2:reset_n, dcc_data_30:reset_n, dcc_data_31:reset_n, dcc_data_3:reset_n, dcc_data_4:reset_n, dcc_data_5:reset_n, dcc_data_6:reset_n, dcc_data_7:reset_n, dcc_data_8:reset_n, dcc_data_9:reset_n, dcc_time_out:reset_n, hps_read_bit:reset_n, jtag_uart:rst_n, ledr:reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, pps_count_out:reset_n, rst_translator:in_reset, sw:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [irq_mapper_002:reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	soc_system_dcc_data_0 dcc_data_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_0_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_0_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_1 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_1_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_1_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_10 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_10_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_10_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_10_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_10_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_10_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_10_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver12_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_11 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_11_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_11_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_11_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_11_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_11_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_11_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver13_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_12 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_12_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_12_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_12_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_12_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_12_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_12_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver14_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_13 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_13_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_13_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_13_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_13_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_13_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_13_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver15_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_14 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_14_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_14_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_14_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_14_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_14_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_14_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver16_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_15 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_15_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_15_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_15_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_15_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_15_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_15_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver17_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_16 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_16_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_16_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_16_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_16_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_16_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_16_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver15_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_17 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_17_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_17_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_17_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_17_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_17_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_17_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver0_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_18 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_18_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_18_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_18_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_18_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_18_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_18_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver1_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_19 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_19_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_19_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_19_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_19_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_19_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_19_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver2_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_2 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_2_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_2_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_20 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_20_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_20_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_20_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_20_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_20_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_20_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver3_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_21 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_21_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_21_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_21_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_21_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_21_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_21_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver4_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_22 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_22_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_22_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_22_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_22_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_22_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_22_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver5_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_23 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_23_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_23_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_23_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_23_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_23_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_23_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver6_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_24 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_24_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_24_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_24_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_24_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_24_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_24_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver7_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_25 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_25_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_25_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_25_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_25_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_25_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_25_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver8_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_26 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_26_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_26_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_26_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_26_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_26_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_26_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver9_irq)                 //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_27 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_27_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_27_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_27_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_27_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_27_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_27_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver10_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_28 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_28_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_28_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_28_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_28_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_28_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_28_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver11_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_29 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_29_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_29_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_29_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_29_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_29_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_29_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver12_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_3 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_3_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_3_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_30 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_30_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_30_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_30_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_30_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_30_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_30_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver13_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_31 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_31_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_31_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_31_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_31_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_31_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_31_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_001_receiver14_irq)                //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_4 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_4_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_4_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_5 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_5_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_5_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver7_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_6 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_6_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_6_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver8_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_7 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_7_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_7_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver9_irq)                    //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_8 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_8_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_8_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver10_irq)                   //                 irq.irq
	);

	soc_system_dcc_data_0 dcc_data_9 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_dcc_data_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_data_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_data_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_data_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_data_9_s1_readdata),   //                    .readdata
		.in_port    (dcc_data_9_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver11_irq)                   //                 irq.irq
	);

	soc_system_dcc_time_out dcc_time_out (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_dcc_time_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dcc_time_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dcc_time_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dcc_time_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dcc_time_out_s1_readdata),   //                    .readdata
		.in_port    (dcc_time_out_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                      //                 irq.irq
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),      //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),     // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),      //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),  //   f2h_stm_hw_events.stm_hwevents
		.f2h_dma_req0_req         (hps_0_f2h_dma_req0_dma_req),            //        f2h_dma_req0.dma_req
		.f2h_dma_req0_single      (hps_0_f2h_dma_req0_dma_single),         //                    .dma_single
		.f2h_dma_req0_ack         (hps_0_f2h_dma_req0_dma_ack),            //                    .dma_ack
		.f2h_dma_req1_req         (hps_0_f2h_dma_req1_dma_req),            //        f2h_dma_req1.dma_req
		.f2h_dma_req1_single      (hps_0_f2h_dma_req1_dma_single),         //                    .dma_single
		.f2h_dma_req1_ack         (hps_0_f2h_dma_req1_dma_ack),            //                    .dma_ack
		.mem_a                    (memory_mem_a),                          //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                         //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                         //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                       //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                        //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                       //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                      //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                      //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                       //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                    //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                         //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                        //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                      //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                        //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                         //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                      //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK), //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),   //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),   //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),   //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),   //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),   //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),   //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),    //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL), //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL), //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK), //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),   //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),   //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),   //                    .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),     //                    .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),     //                    .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),     //                    .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),     //                    .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),     //                    .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),     //                    .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),     //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),      //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),      //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),     //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),      //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),      //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),      //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),      //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),      //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),      //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),      //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),      //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),      //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),      //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),     //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),     //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),     //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),     //                    .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_0_hps_io_hps_io_spim0_inst_CLK),    //                    .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_0_hps_io_hps_io_spim0_inst_MOSI),   //                    .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_0_hps_io_hps_io_spim0_inst_MISO),   //                    .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_0_hps_io_hps_io_spim0_inst_SS0),    //                    .hps_io_spim0_inst_SS0
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),    //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),   //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),   //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),    //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),     //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),     //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),     //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),     //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),     //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),     //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),  //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),  //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO37  (hps_0_hps_io_hps_io_gpio_inst_GPIO37),  //                    .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),  //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),  //                    .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO44  (hps_0_hps_io_hps_io_gpio_inst_GPIO44),  //                    .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),  //                    .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),  //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),  //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),  //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),               //           h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                               //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                                      //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                                      //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (),                                      //                    .waitrequest
		.f2h_sdram0_READDATA      (),                                      //                    .readdata
		.f2h_sdram0_READDATAVALID (),                                      //                    .readdatavalid
		.f2h_sdram0_READ          (),                                      //                    .read
		.f2h_sdram0_WRITEDATA     (),                                      //                    .writedata
		.f2h_sdram0_BYTEENABLE    (),                                      //                    .byteenable
		.f2h_sdram0_WRITE         (),                                      //                    .write
		.h2f_axi_clk              (clk_clk),                               //       h2f_axi_clock.clk
		.h2f_AWID                 (),                                      //      h2f_axi_master.awid
		.h2f_AWADDR               (),                                      //                    .awaddr
		.h2f_AWLEN                (),                                      //                    .awlen
		.h2f_AWSIZE               (),                                      //                    .awsize
		.h2f_AWBURST              (),                                      //                    .awburst
		.h2f_AWLOCK               (),                                      //                    .awlock
		.h2f_AWCACHE              (),                                      //                    .awcache
		.h2f_AWPROT               (),                                      //                    .awprot
		.h2f_AWVALID              (),                                      //                    .awvalid
		.h2f_AWREADY              (),                                      //                    .awready
		.h2f_WID                  (),                                      //                    .wid
		.h2f_WDATA                (),                                      //                    .wdata
		.h2f_WSTRB                (),                                      //                    .wstrb
		.h2f_WLAST                (),                                      //                    .wlast
		.h2f_WVALID               (),                                      //                    .wvalid
		.h2f_WREADY               (),                                      //                    .wready
		.h2f_BID                  (),                                      //                    .bid
		.h2f_BRESP                (),                                      //                    .bresp
		.h2f_BVALID               (),                                      //                    .bvalid
		.h2f_BREADY               (),                                      //                    .bready
		.h2f_ARID                 (),                                      //                    .arid
		.h2f_ARADDR               (),                                      //                    .araddr
		.h2f_ARLEN                (),                                      //                    .arlen
		.h2f_ARSIZE               (),                                      //                    .arsize
		.h2f_ARBURST              (),                                      //                    .arburst
		.h2f_ARLOCK               (),                                      //                    .arlock
		.h2f_ARCACHE              (),                                      //                    .arcache
		.h2f_ARPROT               (),                                      //                    .arprot
		.h2f_ARVALID              (),                                      //                    .arvalid
		.h2f_ARREADY              (),                                      //                    .arready
		.h2f_RID                  (),                                      //                    .rid
		.h2f_RDATA                (),                                      //                    .rdata
		.h2f_RRESP                (),                                      //                    .rresp
		.h2f_RLAST                (),                                      //                    .rlast
		.h2f_RVALID               (),                                      //                    .rvalid
		.h2f_RREADY               (),                                      //                    .rready
		.f2h_axi_clk              (clk_clk),                               //       f2h_axi_clock.clk
		.f2h_AWID                 (),                                      //       f2h_axi_slave.awid
		.f2h_AWADDR               (),                                      //                    .awaddr
		.f2h_AWLEN                (),                                      //                    .awlen
		.f2h_AWSIZE               (),                                      //                    .awsize
		.f2h_AWBURST              (),                                      //                    .awburst
		.f2h_AWLOCK               (),                                      //                    .awlock
		.f2h_AWCACHE              (),                                      //                    .awcache
		.f2h_AWPROT               (),                                      //                    .awprot
		.f2h_AWVALID              (),                                      //                    .awvalid
		.f2h_AWREADY              (),                                      //                    .awready
		.f2h_AWUSER               (),                                      //                    .awuser
		.f2h_WID                  (),                                      //                    .wid
		.f2h_WDATA                (),                                      //                    .wdata
		.f2h_WSTRB                (),                                      //                    .wstrb
		.f2h_WLAST                (),                                      //                    .wlast
		.f2h_WVALID               (),                                      //                    .wvalid
		.f2h_WREADY               (),                                      //                    .wready
		.f2h_BID                  (),                                      //                    .bid
		.f2h_BRESP                (),                                      //                    .bresp
		.f2h_BVALID               (),                                      //                    .bvalid
		.f2h_BREADY               (),                                      //                    .bready
		.f2h_ARID                 (),                                      //                    .arid
		.f2h_ARADDR               (),                                      //                    .araddr
		.f2h_ARLEN                (),                                      //                    .arlen
		.f2h_ARSIZE               (),                                      //                    .arsize
		.f2h_ARBURST              (),                                      //                    .arburst
		.f2h_ARLOCK               (),                                      //                    .arlock
		.f2h_ARCACHE              (),                                      //                    .arcache
		.f2h_ARPROT               (),                                      //                    .arprot
		.f2h_ARVALID              (),                                      //                    .arvalid
		.f2h_ARREADY              (),                                      //                    .arready
		.f2h_ARUSER               (),                                      //                    .aruser
		.f2h_RID                  (),                                      //                    .rid
		.f2h_RDATA                (),                                      //                    .rdata
		.f2h_RRESP                (),                                      //                    .rresp
		.f2h_RLAST                (),                                      //                    .rlast
		.f2h_RVALID               (),                                      //                    .rvalid
		.f2h_RREADY               (),                                      //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                               //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),          //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),        //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),         //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),        //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),       //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),        //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),       //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),        //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),       //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),       //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),           //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),         //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),         //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),         //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),        //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),        //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),           //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),         //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),        //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),        //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),          //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),        //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),         //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),        //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),       //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),        //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),       //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),        //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),       //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),       //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),           //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),         //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),         //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),         //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),        //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),        //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                    //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                     //            f2h_irq1.irq
	);

	soc_system_hps_read_bit hps_read_bit (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_hps_read_bit_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hps_read_bit_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hps_read_bit_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hps_read_bit_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hps_read_bit_s1_readdata),   //                    .readdata
		.out_port   (hps_read_bit_external_connection_export)       // external_connection.export
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                               //               irq.irq
	);

	soc_system_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	soc_system_nios2_gen2 nios2_gen2 (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	soc_system_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	soc_system_dcc_data_0 pps_count_out (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pps_count_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pps_count_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pps_count_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pps_count_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pps_count_out_s1_readdata),   //                    .readdata
		.in_port    (pps_count_out_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver18_irq)                      //                 irq.irq
	);

	soc_system_sw sw (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver0_irq)            //                 irq.irq
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver0_irq)           //   irq.irq
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                (clk_clk),                                                   //                              clk_50_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                        //  nios2_gen2_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                    //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                 //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                 //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                       //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                   //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                              //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                      //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                  //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                //                                        .debugaccess
		.nios2_gen2_data_master_address                (nios2_gen2_data_master_address),                            //                  nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest            (nios2_gen2_data_master_waitrequest),                        //                                        .waitrequest
		.nios2_gen2_data_master_byteenable             (nios2_gen2_data_master_byteenable),                         //                                        .byteenable
		.nios2_gen2_data_master_read                   (nios2_gen2_data_master_read),                               //                                        .read
		.nios2_gen2_data_master_readdata               (nios2_gen2_data_master_readdata),                           //                                        .readdata
		.nios2_gen2_data_master_write                  (nios2_gen2_data_master_write),                              //                                        .write
		.nios2_gen2_data_master_writedata              (nios2_gen2_data_master_writedata),                          //                                        .writedata
		.nios2_gen2_data_master_debugaccess            (nios2_gen2_data_master_debugaccess),                        //                                        .debugaccess
		.nios2_gen2_instruction_master_address         (nios2_gen2_instruction_master_address),                     //           nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest     (nios2_gen2_instruction_master_waitrequest),                 //                                        .waitrequest
		.nios2_gen2_instruction_master_read            (nios2_gen2_instruction_master_read),                        //                                        .read
		.nios2_gen2_instruction_master_readdata        (nios2_gen2_instruction_master_readdata),                    //                                        .readdata
		.dcc_data_0_s1_address                         (mm_interconnect_0_dcc_data_0_s1_address),                   //                           dcc_data_0_s1.address
		.dcc_data_0_s1_write                           (mm_interconnect_0_dcc_data_0_s1_write),                     //                                        .write
		.dcc_data_0_s1_readdata                        (mm_interconnect_0_dcc_data_0_s1_readdata),                  //                                        .readdata
		.dcc_data_0_s1_writedata                       (mm_interconnect_0_dcc_data_0_s1_writedata),                 //                                        .writedata
		.dcc_data_0_s1_chipselect                      (mm_interconnect_0_dcc_data_0_s1_chipselect),                //                                        .chipselect
		.dcc_data_1_s1_address                         (mm_interconnect_0_dcc_data_1_s1_address),                   //                           dcc_data_1_s1.address
		.dcc_data_1_s1_write                           (mm_interconnect_0_dcc_data_1_s1_write),                     //                                        .write
		.dcc_data_1_s1_readdata                        (mm_interconnect_0_dcc_data_1_s1_readdata),                  //                                        .readdata
		.dcc_data_1_s1_writedata                       (mm_interconnect_0_dcc_data_1_s1_writedata),                 //                                        .writedata
		.dcc_data_1_s1_chipselect                      (mm_interconnect_0_dcc_data_1_s1_chipselect),                //                                        .chipselect
		.dcc_data_10_s1_address                        (mm_interconnect_0_dcc_data_10_s1_address),                  //                          dcc_data_10_s1.address
		.dcc_data_10_s1_write                          (mm_interconnect_0_dcc_data_10_s1_write),                    //                                        .write
		.dcc_data_10_s1_readdata                       (mm_interconnect_0_dcc_data_10_s1_readdata),                 //                                        .readdata
		.dcc_data_10_s1_writedata                      (mm_interconnect_0_dcc_data_10_s1_writedata),                //                                        .writedata
		.dcc_data_10_s1_chipselect                     (mm_interconnect_0_dcc_data_10_s1_chipselect),               //                                        .chipselect
		.dcc_data_11_s1_address                        (mm_interconnect_0_dcc_data_11_s1_address),                  //                          dcc_data_11_s1.address
		.dcc_data_11_s1_write                          (mm_interconnect_0_dcc_data_11_s1_write),                    //                                        .write
		.dcc_data_11_s1_readdata                       (mm_interconnect_0_dcc_data_11_s1_readdata),                 //                                        .readdata
		.dcc_data_11_s1_writedata                      (mm_interconnect_0_dcc_data_11_s1_writedata),                //                                        .writedata
		.dcc_data_11_s1_chipselect                     (mm_interconnect_0_dcc_data_11_s1_chipselect),               //                                        .chipselect
		.dcc_data_12_s1_address                        (mm_interconnect_0_dcc_data_12_s1_address),                  //                          dcc_data_12_s1.address
		.dcc_data_12_s1_write                          (mm_interconnect_0_dcc_data_12_s1_write),                    //                                        .write
		.dcc_data_12_s1_readdata                       (mm_interconnect_0_dcc_data_12_s1_readdata),                 //                                        .readdata
		.dcc_data_12_s1_writedata                      (mm_interconnect_0_dcc_data_12_s1_writedata),                //                                        .writedata
		.dcc_data_12_s1_chipselect                     (mm_interconnect_0_dcc_data_12_s1_chipselect),               //                                        .chipselect
		.dcc_data_13_s1_address                        (mm_interconnect_0_dcc_data_13_s1_address),                  //                          dcc_data_13_s1.address
		.dcc_data_13_s1_write                          (mm_interconnect_0_dcc_data_13_s1_write),                    //                                        .write
		.dcc_data_13_s1_readdata                       (mm_interconnect_0_dcc_data_13_s1_readdata),                 //                                        .readdata
		.dcc_data_13_s1_writedata                      (mm_interconnect_0_dcc_data_13_s1_writedata),                //                                        .writedata
		.dcc_data_13_s1_chipselect                     (mm_interconnect_0_dcc_data_13_s1_chipselect),               //                                        .chipselect
		.dcc_data_14_s1_address                        (mm_interconnect_0_dcc_data_14_s1_address),                  //                          dcc_data_14_s1.address
		.dcc_data_14_s1_write                          (mm_interconnect_0_dcc_data_14_s1_write),                    //                                        .write
		.dcc_data_14_s1_readdata                       (mm_interconnect_0_dcc_data_14_s1_readdata),                 //                                        .readdata
		.dcc_data_14_s1_writedata                      (mm_interconnect_0_dcc_data_14_s1_writedata),                //                                        .writedata
		.dcc_data_14_s1_chipselect                     (mm_interconnect_0_dcc_data_14_s1_chipselect),               //                                        .chipselect
		.dcc_data_15_s1_address                        (mm_interconnect_0_dcc_data_15_s1_address),                  //                          dcc_data_15_s1.address
		.dcc_data_15_s1_write                          (mm_interconnect_0_dcc_data_15_s1_write),                    //                                        .write
		.dcc_data_15_s1_readdata                       (mm_interconnect_0_dcc_data_15_s1_readdata),                 //                                        .readdata
		.dcc_data_15_s1_writedata                      (mm_interconnect_0_dcc_data_15_s1_writedata),                //                                        .writedata
		.dcc_data_15_s1_chipselect                     (mm_interconnect_0_dcc_data_15_s1_chipselect),               //                                        .chipselect
		.dcc_data_16_s1_address                        (mm_interconnect_0_dcc_data_16_s1_address),                  //                          dcc_data_16_s1.address
		.dcc_data_16_s1_write                          (mm_interconnect_0_dcc_data_16_s1_write),                    //                                        .write
		.dcc_data_16_s1_readdata                       (mm_interconnect_0_dcc_data_16_s1_readdata),                 //                                        .readdata
		.dcc_data_16_s1_writedata                      (mm_interconnect_0_dcc_data_16_s1_writedata),                //                                        .writedata
		.dcc_data_16_s1_chipselect                     (mm_interconnect_0_dcc_data_16_s1_chipselect),               //                                        .chipselect
		.dcc_data_17_s1_address                        (mm_interconnect_0_dcc_data_17_s1_address),                  //                          dcc_data_17_s1.address
		.dcc_data_17_s1_write                          (mm_interconnect_0_dcc_data_17_s1_write),                    //                                        .write
		.dcc_data_17_s1_readdata                       (mm_interconnect_0_dcc_data_17_s1_readdata),                 //                                        .readdata
		.dcc_data_17_s1_writedata                      (mm_interconnect_0_dcc_data_17_s1_writedata),                //                                        .writedata
		.dcc_data_17_s1_chipselect                     (mm_interconnect_0_dcc_data_17_s1_chipselect),               //                                        .chipselect
		.dcc_data_18_s1_address                        (mm_interconnect_0_dcc_data_18_s1_address),                  //                          dcc_data_18_s1.address
		.dcc_data_18_s1_write                          (mm_interconnect_0_dcc_data_18_s1_write),                    //                                        .write
		.dcc_data_18_s1_readdata                       (mm_interconnect_0_dcc_data_18_s1_readdata),                 //                                        .readdata
		.dcc_data_18_s1_writedata                      (mm_interconnect_0_dcc_data_18_s1_writedata),                //                                        .writedata
		.dcc_data_18_s1_chipselect                     (mm_interconnect_0_dcc_data_18_s1_chipselect),               //                                        .chipselect
		.dcc_data_19_s1_address                        (mm_interconnect_0_dcc_data_19_s1_address),                  //                          dcc_data_19_s1.address
		.dcc_data_19_s1_write                          (mm_interconnect_0_dcc_data_19_s1_write),                    //                                        .write
		.dcc_data_19_s1_readdata                       (mm_interconnect_0_dcc_data_19_s1_readdata),                 //                                        .readdata
		.dcc_data_19_s1_writedata                      (mm_interconnect_0_dcc_data_19_s1_writedata),                //                                        .writedata
		.dcc_data_19_s1_chipselect                     (mm_interconnect_0_dcc_data_19_s1_chipselect),               //                                        .chipselect
		.dcc_data_2_s1_address                         (mm_interconnect_0_dcc_data_2_s1_address),                   //                           dcc_data_2_s1.address
		.dcc_data_2_s1_write                           (mm_interconnect_0_dcc_data_2_s1_write),                     //                                        .write
		.dcc_data_2_s1_readdata                        (mm_interconnect_0_dcc_data_2_s1_readdata),                  //                                        .readdata
		.dcc_data_2_s1_writedata                       (mm_interconnect_0_dcc_data_2_s1_writedata),                 //                                        .writedata
		.dcc_data_2_s1_chipselect                      (mm_interconnect_0_dcc_data_2_s1_chipselect),                //                                        .chipselect
		.dcc_data_20_s1_address                        (mm_interconnect_0_dcc_data_20_s1_address),                  //                          dcc_data_20_s1.address
		.dcc_data_20_s1_write                          (mm_interconnect_0_dcc_data_20_s1_write),                    //                                        .write
		.dcc_data_20_s1_readdata                       (mm_interconnect_0_dcc_data_20_s1_readdata),                 //                                        .readdata
		.dcc_data_20_s1_writedata                      (mm_interconnect_0_dcc_data_20_s1_writedata),                //                                        .writedata
		.dcc_data_20_s1_chipselect                     (mm_interconnect_0_dcc_data_20_s1_chipselect),               //                                        .chipselect
		.dcc_data_21_s1_address                        (mm_interconnect_0_dcc_data_21_s1_address),                  //                          dcc_data_21_s1.address
		.dcc_data_21_s1_write                          (mm_interconnect_0_dcc_data_21_s1_write),                    //                                        .write
		.dcc_data_21_s1_readdata                       (mm_interconnect_0_dcc_data_21_s1_readdata),                 //                                        .readdata
		.dcc_data_21_s1_writedata                      (mm_interconnect_0_dcc_data_21_s1_writedata),                //                                        .writedata
		.dcc_data_21_s1_chipselect                     (mm_interconnect_0_dcc_data_21_s1_chipselect),               //                                        .chipselect
		.dcc_data_22_s1_address                        (mm_interconnect_0_dcc_data_22_s1_address),                  //                          dcc_data_22_s1.address
		.dcc_data_22_s1_write                          (mm_interconnect_0_dcc_data_22_s1_write),                    //                                        .write
		.dcc_data_22_s1_readdata                       (mm_interconnect_0_dcc_data_22_s1_readdata),                 //                                        .readdata
		.dcc_data_22_s1_writedata                      (mm_interconnect_0_dcc_data_22_s1_writedata),                //                                        .writedata
		.dcc_data_22_s1_chipselect                     (mm_interconnect_0_dcc_data_22_s1_chipselect),               //                                        .chipselect
		.dcc_data_23_s1_address                        (mm_interconnect_0_dcc_data_23_s1_address),                  //                          dcc_data_23_s1.address
		.dcc_data_23_s1_write                          (mm_interconnect_0_dcc_data_23_s1_write),                    //                                        .write
		.dcc_data_23_s1_readdata                       (mm_interconnect_0_dcc_data_23_s1_readdata),                 //                                        .readdata
		.dcc_data_23_s1_writedata                      (mm_interconnect_0_dcc_data_23_s1_writedata),                //                                        .writedata
		.dcc_data_23_s1_chipselect                     (mm_interconnect_0_dcc_data_23_s1_chipselect),               //                                        .chipselect
		.dcc_data_24_s1_address                        (mm_interconnect_0_dcc_data_24_s1_address),                  //                          dcc_data_24_s1.address
		.dcc_data_24_s1_write                          (mm_interconnect_0_dcc_data_24_s1_write),                    //                                        .write
		.dcc_data_24_s1_readdata                       (mm_interconnect_0_dcc_data_24_s1_readdata),                 //                                        .readdata
		.dcc_data_24_s1_writedata                      (mm_interconnect_0_dcc_data_24_s1_writedata),                //                                        .writedata
		.dcc_data_24_s1_chipselect                     (mm_interconnect_0_dcc_data_24_s1_chipselect),               //                                        .chipselect
		.dcc_data_25_s1_address                        (mm_interconnect_0_dcc_data_25_s1_address),                  //                          dcc_data_25_s1.address
		.dcc_data_25_s1_write                          (mm_interconnect_0_dcc_data_25_s1_write),                    //                                        .write
		.dcc_data_25_s1_readdata                       (mm_interconnect_0_dcc_data_25_s1_readdata),                 //                                        .readdata
		.dcc_data_25_s1_writedata                      (mm_interconnect_0_dcc_data_25_s1_writedata),                //                                        .writedata
		.dcc_data_25_s1_chipselect                     (mm_interconnect_0_dcc_data_25_s1_chipselect),               //                                        .chipselect
		.dcc_data_26_s1_address                        (mm_interconnect_0_dcc_data_26_s1_address),                  //                          dcc_data_26_s1.address
		.dcc_data_26_s1_write                          (mm_interconnect_0_dcc_data_26_s1_write),                    //                                        .write
		.dcc_data_26_s1_readdata                       (mm_interconnect_0_dcc_data_26_s1_readdata),                 //                                        .readdata
		.dcc_data_26_s1_writedata                      (mm_interconnect_0_dcc_data_26_s1_writedata),                //                                        .writedata
		.dcc_data_26_s1_chipselect                     (mm_interconnect_0_dcc_data_26_s1_chipselect),               //                                        .chipselect
		.dcc_data_27_s1_address                        (mm_interconnect_0_dcc_data_27_s1_address),                  //                          dcc_data_27_s1.address
		.dcc_data_27_s1_write                          (mm_interconnect_0_dcc_data_27_s1_write),                    //                                        .write
		.dcc_data_27_s1_readdata                       (mm_interconnect_0_dcc_data_27_s1_readdata),                 //                                        .readdata
		.dcc_data_27_s1_writedata                      (mm_interconnect_0_dcc_data_27_s1_writedata),                //                                        .writedata
		.dcc_data_27_s1_chipselect                     (mm_interconnect_0_dcc_data_27_s1_chipselect),               //                                        .chipselect
		.dcc_data_28_s1_address                        (mm_interconnect_0_dcc_data_28_s1_address),                  //                          dcc_data_28_s1.address
		.dcc_data_28_s1_write                          (mm_interconnect_0_dcc_data_28_s1_write),                    //                                        .write
		.dcc_data_28_s1_readdata                       (mm_interconnect_0_dcc_data_28_s1_readdata),                 //                                        .readdata
		.dcc_data_28_s1_writedata                      (mm_interconnect_0_dcc_data_28_s1_writedata),                //                                        .writedata
		.dcc_data_28_s1_chipselect                     (mm_interconnect_0_dcc_data_28_s1_chipselect),               //                                        .chipselect
		.dcc_data_29_s1_address                        (mm_interconnect_0_dcc_data_29_s1_address),                  //                          dcc_data_29_s1.address
		.dcc_data_29_s1_write                          (mm_interconnect_0_dcc_data_29_s1_write),                    //                                        .write
		.dcc_data_29_s1_readdata                       (mm_interconnect_0_dcc_data_29_s1_readdata),                 //                                        .readdata
		.dcc_data_29_s1_writedata                      (mm_interconnect_0_dcc_data_29_s1_writedata),                //                                        .writedata
		.dcc_data_29_s1_chipselect                     (mm_interconnect_0_dcc_data_29_s1_chipselect),               //                                        .chipselect
		.dcc_data_3_s1_address                         (mm_interconnect_0_dcc_data_3_s1_address),                   //                           dcc_data_3_s1.address
		.dcc_data_3_s1_write                           (mm_interconnect_0_dcc_data_3_s1_write),                     //                                        .write
		.dcc_data_3_s1_readdata                        (mm_interconnect_0_dcc_data_3_s1_readdata),                  //                                        .readdata
		.dcc_data_3_s1_writedata                       (mm_interconnect_0_dcc_data_3_s1_writedata),                 //                                        .writedata
		.dcc_data_3_s1_chipselect                      (mm_interconnect_0_dcc_data_3_s1_chipselect),                //                                        .chipselect
		.dcc_data_30_s1_address                        (mm_interconnect_0_dcc_data_30_s1_address),                  //                          dcc_data_30_s1.address
		.dcc_data_30_s1_write                          (mm_interconnect_0_dcc_data_30_s1_write),                    //                                        .write
		.dcc_data_30_s1_readdata                       (mm_interconnect_0_dcc_data_30_s1_readdata),                 //                                        .readdata
		.dcc_data_30_s1_writedata                      (mm_interconnect_0_dcc_data_30_s1_writedata),                //                                        .writedata
		.dcc_data_30_s1_chipselect                     (mm_interconnect_0_dcc_data_30_s1_chipselect),               //                                        .chipselect
		.dcc_data_31_s1_address                        (mm_interconnect_0_dcc_data_31_s1_address),                  //                          dcc_data_31_s1.address
		.dcc_data_31_s1_write                          (mm_interconnect_0_dcc_data_31_s1_write),                    //                                        .write
		.dcc_data_31_s1_readdata                       (mm_interconnect_0_dcc_data_31_s1_readdata),                 //                                        .readdata
		.dcc_data_31_s1_writedata                      (mm_interconnect_0_dcc_data_31_s1_writedata),                //                                        .writedata
		.dcc_data_31_s1_chipselect                     (mm_interconnect_0_dcc_data_31_s1_chipselect),               //                                        .chipselect
		.dcc_data_4_s1_address                         (mm_interconnect_0_dcc_data_4_s1_address),                   //                           dcc_data_4_s1.address
		.dcc_data_4_s1_write                           (mm_interconnect_0_dcc_data_4_s1_write),                     //                                        .write
		.dcc_data_4_s1_readdata                        (mm_interconnect_0_dcc_data_4_s1_readdata),                  //                                        .readdata
		.dcc_data_4_s1_writedata                       (mm_interconnect_0_dcc_data_4_s1_writedata),                 //                                        .writedata
		.dcc_data_4_s1_chipselect                      (mm_interconnect_0_dcc_data_4_s1_chipselect),                //                                        .chipselect
		.dcc_data_5_s1_address                         (mm_interconnect_0_dcc_data_5_s1_address),                   //                           dcc_data_5_s1.address
		.dcc_data_5_s1_write                           (mm_interconnect_0_dcc_data_5_s1_write),                     //                                        .write
		.dcc_data_5_s1_readdata                        (mm_interconnect_0_dcc_data_5_s1_readdata),                  //                                        .readdata
		.dcc_data_5_s1_writedata                       (mm_interconnect_0_dcc_data_5_s1_writedata),                 //                                        .writedata
		.dcc_data_5_s1_chipselect                      (mm_interconnect_0_dcc_data_5_s1_chipselect),                //                                        .chipselect
		.dcc_data_6_s1_address                         (mm_interconnect_0_dcc_data_6_s1_address),                   //                           dcc_data_6_s1.address
		.dcc_data_6_s1_write                           (mm_interconnect_0_dcc_data_6_s1_write),                     //                                        .write
		.dcc_data_6_s1_readdata                        (mm_interconnect_0_dcc_data_6_s1_readdata),                  //                                        .readdata
		.dcc_data_6_s1_writedata                       (mm_interconnect_0_dcc_data_6_s1_writedata),                 //                                        .writedata
		.dcc_data_6_s1_chipselect                      (mm_interconnect_0_dcc_data_6_s1_chipselect),                //                                        .chipselect
		.dcc_data_7_s1_address                         (mm_interconnect_0_dcc_data_7_s1_address),                   //                           dcc_data_7_s1.address
		.dcc_data_7_s1_write                           (mm_interconnect_0_dcc_data_7_s1_write),                     //                                        .write
		.dcc_data_7_s1_readdata                        (mm_interconnect_0_dcc_data_7_s1_readdata),                  //                                        .readdata
		.dcc_data_7_s1_writedata                       (mm_interconnect_0_dcc_data_7_s1_writedata),                 //                                        .writedata
		.dcc_data_7_s1_chipselect                      (mm_interconnect_0_dcc_data_7_s1_chipselect),                //                                        .chipselect
		.dcc_data_8_s1_address                         (mm_interconnect_0_dcc_data_8_s1_address),                   //                           dcc_data_8_s1.address
		.dcc_data_8_s1_write                           (mm_interconnect_0_dcc_data_8_s1_write),                     //                                        .write
		.dcc_data_8_s1_readdata                        (mm_interconnect_0_dcc_data_8_s1_readdata),                  //                                        .readdata
		.dcc_data_8_s1_writedata                       (mm_interconnect_0_dcc_data_8_s1_writedata),                 //                                        .writedata
		.dcc_data_8_s1_chipselect                      (mm_interconnect_0_dcc_data_8_s1_chipselect),                //                                        .chipselect
		.dcc_data_9_s1_address                         (mm_interconnect_0_dcc_data_9_s1_address),                   //                           dcc_data_9_s1.address
		.dcc_data_9_s1_write                           (mm_interconnect_0_dcc_data_9_s1_write),                     //                                        .write
		.dcc_data_9_s1_readdata                        (mm_interconnect_0_dcc_data_9_s1_readdata),                  //                                        .readdata
		.dcc_data_9_s1_writedata                       (mm_interconnect_0_dcc_data_9_s1_writedata),                 //                                        .writedata
		.dcc_data_9_s1_chipselect                      (mm_interconnect_0_dcc_data_9_s1_chipselect),                //                                        .chipselect
		.dcc_time_out_s1_address                       (mm_interconnect_0_dcc_time_out_s1_address),                 //                         dcc_time_out_s1.address
		.dcc_time_out_s1_write                         (mm_interconnect_0_dcc_time_out_s1_write),                   //                                        .write
		.dcc_time_out_s1_readdata                      (mm_interconnect_0_dcc_time_out_s1_readdata),                //                                        .readdata
		.dcc_time_out_s1_writedata                     (mm_interconnect_0_dcc_time_out_s1_writedata),               //                                        .writedata
		.dcc_time_out_s1_chipselect                    (mm_interconnect_0_dcc_time_out_s1_chipselect),              //                                        .chipselect
		.hps_read_bit_s1_address                       (mm_interconnect_0_hps_read_bit_s1_address),                 //                         hps_read_bit_s1.address
		.hps_read_bit_s1_write                         (mm_interconnect_0_hps_read_bit_s1_write),                   //                                        .write
		.hps_read_bit_s1_readdata                      (mm_interconnect_0_hps_read_bit_s1_readdata),                //                                        .readdata
		.hps_read_bit_s1_writedata                     (mm_interconnect_0_hps_read_bit_s1_writedata),               //                                        .writedata
		.hps_read_bit_s1_chipselect                    (mm_interconnect_0_hps_read_bit_s1_chipselect),              //                                        .chipselect
		.jtag_uart_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.ledr_s1_address                               (mm_interconnect_0_ledr_s1_address),                         //                                 ledr_s1.address
		.ledr_s1_write                                 (mm_interconnect_0_ledr_s1_write),                           //                                        .write
		.ledr_s1_readdata                              (mm_interconnect_0_ledr_s1_readdata),                        //                                        .readdata
		.ledr_s1_writedata                             (mm_interconnect_0_ledr_s1_writedata),                       //                                        .writedata
		.ledr_s1_chipselect                            (mm_interconnect_0_ledr_s1_chipselect),                      //                                        .chipselect
		.nios2_gen2_debug_mem_slave_address            (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //              nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write              (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                        .write
		.nios2_gen2_debug_mem_slave_read               (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                        .read
		.nios2_gen2_debug_mem_slave_readdata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                        .readdata
		.nios2_gen2_debug_mem_slave_writedata          (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                        .writedata
		.nios2_gen2_debug_mem_slave_byteenable         (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                        .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest        (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                        .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess        (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                        .debugaccess
		.onchip_memory2_s1_address                     (mm_interconnect_0_onchip_memory2_s1_address),               //                       onchip_memory2_s1.address
		.onchip_memory2_s1_write                       (mm_interconnect_0_onchip_memory2_s1_write),                 //                                        .write
		.onchip_memory2_s1_readdata                    (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                        .readdata
		.onchip_memory2_s1_writedata                   (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                        .writedata
		.onchip_memory2_s1_byteenable                  (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                        .byteenable
		.onchip_memory2_s1_chipselect                  (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                        .chipselect
		.onchip_memory2_s1_clken                       (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                        .clken
		.pps_count_out_s1_address                      (mm_interconnect_0_pps_count_out_s1_address),                //                        pps_count_out_s1.address
		.pps_count_out_s1_write                        (mm_interconnect_0_pps_count_out_s1_write),                  //                                        .write
		.pps_count_out_s1_readdata                     (mm_interconnect_0_pps_count_out_s1_readdata),               //                                        .readdata
		.pps_count_out_s1_writedata                    (mm_interconnect_0_pps_count_out_s1_writedata),              //                                        .writedata
		.pps_count_out_s1_chipselect                   (mm_interconnect_0_pps_count_out_s1_chipselect),             //                                        .chipselect
		.sw_s1_address                                 (mm_interconnect_0_sw_s1_address),                           //                                   sw_s1.address
		.sw_s1_write                                   (mm_interconnect_0_sw_s1_write),                             //                                        .write
		.sw_s1_readdata                                (mm_interconnect_0_sw_s1_readdata),                          //                                        .readdata
		.sw_s1_writedata                               (mm_interconnect_0_sw_s1_writedata),                         //                                        .writedata
		.sw_s1_chipselect                              (mm_interconnect_0_sw_s1_chipselect),                        //                                        .chipselect
		.sysid_qsys_control_slave_address              (mm_interconnect_0_sysid_qsys_control_slave_address),        //                sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata             (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                        .readdata
		.timer_s1_address                              (mm_interconnect_0_timer_s1_address),                        //                                timer_s1.address
		.timer_s1_write                                (mm_interconnect_0_timer_s1_write),                          //                                        .write
		.timer_s1_readdata                             (mm_interconnect_0_timer_s1_readdata),                       //                                        .readdata
		.timer_s1_writedata                            (mm_interconnect_0_timer_s1_writedata),                      //                                        .writedata
		.timer_s1_chipselect                           (mm_interconnect_0_timer_s1_chipselect)                      //                                        .chipselect
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                   //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                 //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                  //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                 //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                 //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                 //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                    //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                  //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                  //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                  //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                 //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                 //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                    //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                  //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                 //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                 //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                   //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                 //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                  //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                 //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                 //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                 //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                    //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                  //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                  //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                  //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                 //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                 //                                                              .rready
		.clk_50_clk_clk                                                      (clk_clk),                                        //                                                    clk_50_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),             // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset                       (rst_controller_reset_out_reset),                 //                       mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_s0_address                                              (mm_interconnect_1_mm_bridge_0_s0_address),       //                                                mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                                (mm_interconnect_1_mm_bridge_0_s0_write),         //                                                              .write
		.mm_bridge_0_s0_read                                                 (mm_interconnect_1_mm_bridge_0_s0_read),          //                                                              .read
		.mm_bridge_0_s0_readdata                                             (mm_interconnect_1_mm_bridge_0_s0_readdata),      //                                                              .readdata
		.mm_bridge_0_s0_writedata                                            (mm_interconnect_1_mm_bridge_0_s0_writedata),     //                                                              .writedata
		.mm_bridge_0_s0_burstcount                                           (mm_interconnect_1_mm_bridge_0_s0_burstcount),    //                                                              .burstcount
		.mm_bridge_0_s0_byteenable                                           (mm_interconnect_1_mm_bridge_0_s0_byteenable),    //                                                              .byteenable
		.mm_bridge_0_s0_readdatavalid                                        (mm_interconnect_1_mm_bridge_0_s0_readdatavalid), //                                                              .readdatavalid
		.mm_bridge_0_s0_waitrequest                                          (mm_interconnect_1_mm_bridge_0_s0_waitrequest),   //                                                              .waitrequest
		.mm_bridge_0_s0_debugaccess                                          (mm_interconnect_1_mm_bridge_0_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_irq_mapper irq_mapper (
		.clk            (),                          //        clk.clk
		.reset          (),                          //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),  //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),  //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),  //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),  //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),  //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),  //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),  //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),  //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),  //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),  //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq), // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq), // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq), // receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq), // receiver13.irq
		.receiver14_irq (irq_mapper_receiver14_irq), // receiver14.irq
		.receiver15_irq (irq_mapper_receiver15_irq), // receiver15.irq
		.receiver16_irq (irq_mapper_receiver16_irq), // receiver16.irq
		.receiver17_irq (irq_mapper_receiver17_irq), // receiver17.irq
		.receiver18_irq (irq_mapper_receiver18_irq), // receiver18.irq
		.sender_irq     (hps_0_f2h_irq0_irq)         //     sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk            (),                              //        clk.clk
		.reset          (),                              //  clk_reset.reset
		.receiver0_irq  (irq_mapper_001_receiver0_irq),  //  receiver0.irq
		.receiver1_irq  (irq_mapper_001_receiver1_irq),  //  receiver1.irq
		.receiver2_irq  (irq_mapper_001_receiver2_irq),  //  receiver2.irq
		.receiver3_irq  (irq_mapper_001_receiver3_irq),  //  receiver3.irq
		.receiver4_irq  (irq_mapper_001_receiver4_irq),  //  receiver4.irq
		.receiver5_irq  (irq_mapper_001_receiver5_irq),  //  receiver5.irq
		.receiver6_irq  (irq_mapper_001_receiver6_irq),  //  receiver6.irq
		.receiver7_irq  (irq_mapper_001_receiver7_irq),  //  receiver7.irq
		.receiver8_irq  (irq_mapper_001_receiver8_irq),  //  receiver8.irq
		.receiver9_irq  (irq_mapper_001_receiver9_irq),  //  receiver9.irq
		.receiver10_irq (irq_mapper_001_receiver10_irq), // receiver10.irq
		.receiver11_irq (irq_mapper_001_receiver11_irq), // receiver11.irq
		.receiver12_irq (irq_mapper_001_receiver12_irq), // receiver12.irq
		.receiver13_irq (irq_mapper_001_receiver13_irq), // receiver13.irq
		.receiver14_irq (irq_mapper_001_receiver14_irq), // receiver14.irq
		.receiver15_irq (irq_mapper_001_receiver15_irq), // receiver15.irq
		.sender_irq     (hps_0_f2h_irq1_irq)             //     sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_debug_reset_request_reset),   // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
