// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: Shift.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Shift (
	aclr,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps10x,
	taps11x,
	taps12x,
	taps13x,
	taps14x,
	taps15x,
	taps16x,
	taps17x,
	taps18x,
	taps19x,
	taps1x,
	taps20x,
	taps21x,
	taps22x,
	taps23x,
	taps24x,
	taps25x,
	taps26x,
	taps27x,
	taps28x,
	taps29x,
	taps2x,
	taps30x,
	taps31x,
	taps32x,
	taps33x,
	taps34x,
	taps35x,
	taps36x,
	taps37x,
	taps38x,
	taps39x,
	taps3x,
	taps40x,
	taps41x,
	taps42x,
	taps43x,
	taps44x,
	taps45x,
	taps46x,
	taps47x,
	taps48x,
	taps49x,
	taps4x,
	taps50x,
	taps51x,
	taps52x,
	taps53x,
	taps54x,
	taps55x,
	taps56x,
	taps57x,
	taps58x,
	taps59x,
	taps5x,
	taps60x,
	taps61x,
	taps62x,
	taps63x,
	taps64x,
	taps65x,
	taps66x,
	taps67x,
	taps68x,
	taps69x,
	taps6x,
	taps70x,
	taps71x,
	taps72x,
	taps73x,
	taps74x,
	taps75x,
	taps76x,
	taps77x,
	taps78x,
	taps79x,
	taps7x,
	taps80x,
	taps81x,
	taps82x,
	taps83x,
	taps84x,
	taps85x,
	taps86x,
	taps87x,
	taps88x,
	taps89x,
	taps8x,
	taps90x,
	taps91x,
	taps92x,
	taps93x,
	taps94x,
	taps95x,
	taps9x);

	input	  aclr;
	input	  clock;
	input	[15:0]  shiftin;
	output	[15:0]  shiftout;
	output	[15:0]  taps0x;
	output	[15:0]  taps10x;
	output	[15:0]  taps11x;
	output	[15:0]  taps12x;
	output	[15:0]  taps13x;
	output	[15:0]  taps14x;
	output	[15:0]  taps15x;
	output	[15:0]  taps16x;
	output	[15:0]  taps17x;
	output	[15:0]  taps18x;
	output	[15:0]  taps19x;
	output	[15:0]  taps1x;
	output	[15:0]  taps20x;
	output	[15:0]  taps21x;
	output	[15:0]  taps22x;
	output	[15:0]  taps23x;
	output	[15:0]  taps24x;
	output	[15:0]  taps25x;
	output	[15:0]  taps26x;
	output	[15:0]  taps27x;
	output	[15:0]  taps28x;
	output	[15:0]  taps29x;
	output	[15:0]  taps2x;
	output	[15:0]  taps30x;
	output	[15:0]  taps31x;
	output	[15:0]  taps32x;
	output	[15:0]  taps33x;
	output	[15:0]  taps34x;
	output	[15:0]  taps35x;
	output	[15:0]  taps36x;
	output	[15:0]  taps37x;
	output	[15:0]  taps38x;
	output	[15:0]  taps39x;
	output	[15:0]  taps3x;
	output	[15:0]  taps40x;
	output	[15:0]  taps41x;
	output	[15:0]  taps42x;
	output	[15:0]  taps43x;
	output	[15:0]  taps44x;
	output	[15:0]  taps45x;
	output	[15:0]  taps46x;
	output	[15:0]  taps47x;
	output	[15:0]  taps48x;
	output	[15:0]  taps49x;
	output	[15:0]  taps4x;
	output	[15:0]  taps50x;
	output	[15:0]  taps51x;
	output	[15:0]  taps52x;
	output	[15:0]  taps53x;
	output	[15:0]  taps54x;
	output	[15:0]  taps55x;
	output	[15:0]  taps56x;
	output	[15:0]  taps57x;
	output	[15:0]  taps58x;
	output	[15:0]  taps59x;
	output	[15:0]  taps5x;
	output	[15:0]  taps60x;
	output	[15:0]  taps61x;
	output	[15:0]  taps62x;
	output	[15:0]  taps63x;
	output	[15:0]  taps64x;
	output	[15:0]  taps65x;
	output	[15:0]  taps66x;
	output	[15:0]  taps67x;
	output	[15:0]  taps68x;
	output	[15:0]  taps69x;
	output	[15:0]  taps6x;
	output	[15:0]  taps70x;
	output	[15:0]  taps71x;
	output	[15:0]  taps72x;
	output	[15:0]  taps73x;
	output	[15:0]  taps74x;
	output	[15:0]  taps75x;
	output	[15:0]  taps76x;
	output	[15:0]  taps77x;
	output	[15:0]  taps78x;
	output	[15:0]  taps79x;
	output	[15:0]  taps7x;
	output	[15:0]  taps80x;
	output	[15:0]  taps81x;
	output	[15:0]  taps82x;
	output	[15:0]  taps83x;
	output	[15:0]  taps84x;
	output	[15:0]  taps85x;
	output	[15:0]  taps86x;
	output	[15:0]  taps87x;
	output	[15:0]  taps88x;
	output	[15:0]  taps89x;
	output	[15:0]  taps8x;
	output	[15:0]  taps90x;
	output	[15:0]  taps91x;
	output	[15:0]  taps92x;
	output	[15:0]  taps93x;
	output	[15:0]  taps94x;
	output	[15:0]  taps95x;
	output	[15:0]  taps9x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  aclr;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [15:0] sub_wire0;
	wire [1535:0] sub_wire1;
	wire [15:0] shiftout = sub_wire0[15:0];
	wire [159:144] sub_wire191 = sub_wire1[159:144];
	wire [1535:1520] sub_wire190 = sub_wire1[1535:1520];
	wire [1535:1520] sub_wire189 = sub_wire190[1535:1520];
	wire [1519:1504] sub_wire188 = sub_wire1[1519:1504];
	wire [1519:1504] sub_wire187 = sub_wire188[1519:1504];
	wire [1503:1488] sub_wire186 = sub_wire1[1503:1488];
	wire [1503:1488] sub_wire185 = sub_wire186[1503:1488];
	wire [1487:1472] sub_wire184 = sub_wire1[1487:1472];
	wire [1487:1472] sub_wire183 = sub_wire184[1487:1472];
	wire [1471:1456] sub_wire182 = sub_wire1[1471:1456];
	wire [1471:1456] sub_wire181 = sub_wire182[1471:1456];
	wire [1455:1440] sub_wire180 = sub_wire1[1455:1440];
	wire [1455:1440] sub_wire179 = sub_wire180[1455:1440];
	wire [143:128] sub_wire178 = sub_wire1[143:128];
	wire [143:128] sub_wire177 = sub_wire178[143:128];
	wire [1439:1424] sub_wire176 = sub_wire1[1439:1424];
	wire [1439:1424] sub_wire175 = sub_wire176[1439:1424];
	wire [1423:1408] sub_wire174 = sub_wire1[1423:1408];
	wire [1423:1408] sub_wire173 = sub_wire174[1423:1408];
	wire [1407:1392] sub_wire172 = sub_wire1[1407:1392];
	wire [1407:1392] sub_wire171 = sub_wire172[1407:1392];
	wire [1391:1376] sub_wire170 = sub_wire1[1391:1376];
	wire [1391:1376] sub_wire169 = sub_wire170[1391:1376];
	wire [1375:1360] sub_wire168 = sub_wire1[1375:1360];
	wire [1375:1360] sub_wire167 = sub_wire168[1375:1360];
	wire [1359:1344] sub_wire166 = sub_wire1[1359:1344];
	wire [1359:1344] sub_wire165 = sub_wire166[1359:1344];
	wire [1343:1328] sub_wire164 = sub_wire1[1343:1328];
	wire [1343:1328] sub_wire163 = sub_wire164[1343:1328];
	wire [1327:1312] sub_wire162 = sub_wire1[1327:1312];
	wire [1327:1312] sub_wire161 = sub_wire162[1327:1312];
	wire [1311:1296] sub_wire160 = sub_wire1[1311:1296];
	wire [1311:1296] sub_wire159 = sub_wire160[1311:1296];
	wire [1295:1280] sub_wire158 = sub_wire1[1295:1280];
	wire [1295:1280] sub_wire157 = sub_wire158[1295:1280];
	wire [127:112] sub_wire156 = sub_wire1[127:112];
	wire [127:112] sub_wire155 = sub_wire156[127:112];
	wire [1279:1264] sub_wire154 = sub_wire1[1279:1264];
	wire [1279:1264] sub_wire153 = sub_wire154[1279:1264];
	wire [1263:1248] sub_wire152 = sub_wire1[1263:1248];
	wire [1263:1248] sub_wire151 = sub_wire152[1263:1248];
	wire [1247:1232] sub_wire150 = sub_wire1[1247:1232];
	wire [1247:1232] sub_wire149 = sub_wire150[1247:1232];
	wire [1231:1216] sub_wire148 = sub_wire1[1231:1216];
	wire [1231:1216] sub_wire147 = sub_wire148[1231:1216];
	wire [1215:1200] sub_wire146 = sub_wire1[1215:1200];
	wire [1215:1200] sub_wire145 = sub_wire146[1215:1200];
	wire [1199:1184] sub_wire144 = sub_wire1[1199:1184];
	wire [1199:1184] sub_wire143 = sub_wire144[1199:1184];
	wire [1183:1168] sub_wire142 = sub_wire1[1183:1168];
	wire [1183:1168] sub_wire141 = sub_wire142[1183:1168];
	wire [1167:1152] sub_wire140 = sub_wire1[1167:1152];
	wire [1167:1152] sub_wire139 = sub_wire140[1167:1152];
	wire [1151:1136] sub_wire138 = sub_wire1[1151:1136];
	wire [1151:1136] sub_wire137 = sub_wire138[1151:1136];
	wire [1135:1120] sub_wire136 = sub_wire1[1135:1120];
	wire [1135:1120] sub_wire135 = sub_wire136[1135:1120];
	wire [111:96] sub_wire134 = sub_wire1[111:96];
	wire [111:96] sub_wire133 = sub_wire134[111:96];
	wire [1119:1104] sub_wire132 = sub_wire1[1119:1104];
	wire [1119:1104] sub_wire131 = sub_wire132[1119:1104];
	wire [1103:1088] sub_wire130 = sub_wire1[1103:1088];
	wire [1103:1088] sub_wire129 = sub_wire130[1103:1088];
	wire [1087:1072] sub_wire128 = sub_wire1[1087:1072];
	wire [1087:1072] sub_wire127 = sub_wire128[1087:1072];
	wire [1071:1056] sub_wire126 = sub_wire1[1071:1056];
	wire [1071:1056] sub_wire125 = sub_wire126[1071:1056];
	wire [1055:1040] sub_wire124 = sub_wire1[1055:1040];
	wire [1055:1040] sub_wire123 = sub_wire124[1055:1040];
	wire [1039:1024] sub_wire122 = sub_wire1[1039:1024];
	wire [1039:1024] sub_wire121 = sub_wire122[1039:1024];
	wire [1023:1008] sub_wire120 = sub_wire1[1023:1008];
	wire [1023:1008] sub_wire119 = sub_wire120[1023:1008];
	wire [1007:992] sub_wire118 = sub_wire1[1007:992];
	wire [1007:992] sub_wire117 = sub_wire118[1007:992];
	wire [991:976] sub_wire116 = sub_wire1[991:976];
	wire [991:976] sub_wire115 = sub_wire116[991:976];
	wire [975:960] sub_wire114 = sub_wire1[975:960];
	wire [975:960] sub_wire113 = sub_wire114[975:960];
	wire [95:80] sub_wire112 = sub_wire1[95:80];
	wire [95:80] sub_wire111 = sub_wire112[95:80];
	wire [959:944] sub_wire110 = sub_wire1[959:944];
	wire [959:944] sub_wire109 = sub_wire110[959:944];
	wire [943:928] sub_wire108 = sub_wire1[943:928];
	wire [943:928] sub_wire107 = sub_wire108[943:928];
	wire [927:912] sub_wire106 = sub_wire1[927:912];
	wire [927:912] sub_wire105 = sub_wire106[927:912];
	wire [911:896] sub_wire104 = sub_wire1[911:896];
	wire [911:896] sub_wire103 = sub_wire104[911:896];
	wire [895:880] sub_wire102 = sub_wire1[895:880];
	wire [895:880] sub_wire101 = sub_wire102[895:880];
	wire [879:864] sub_wire100 = sub_wire1[879:864];
	wire [879:864] sub_wire99 = sub_wire100[879:864];
	wire [863:848] sub_wire98 = sub_wire1[863:848];
	wire [863:848] sub_wire97 = sub_wire98[863:848];
	wire [847:832] sub_wire96 = sub_wire1[847:832];
	wire [847:832] sub_wire95 = sub_wire96[847:832];
	wire [831:816] sub_wire94 = sub_wire1[831:816];
	wire [831:816] sub_wire93 = sub_wire94[831:816];
	wire [815:800] sub_wire92 = sub_wire1[815:800];
	wire [815:800] sub_wire91 = sub_wire92[815:800];
	wire [79:64] sub_wire90 = sub_wire1[79:64];
	wire [79:64] sub_wire89 = sub_wire90[79:64];
	wire [799:784] sub_wire88 = sub_wire1[799:784];
	wire [799:784] sub_wire87 = sub_wire88[799:784];
	wire [783:768] sub_wire86 = sub_wire1[783:768];
	wire [783:768] sub_wire85 = sub_wire86[783:768];
	wire [767:752] sub_wire84 = sub_wire1[767:752];
	wire [767:752] sub_wire83 = sub_wire84[767:752];
	wire [751:736] sub_wire82 = sub_wire1[751:736];
	wire [751:736] sub_wire81 = sub_wire82[751:736];
	wire [735:720] sub_wire80 = sub_wire1[735:720];
	wire [735:720] sub_wire79 = sub_wire80[735:720];
	wire [719:704] sub_wire78 = sub_wire1[719:704];
	wire [719:704] sub_wire77 = sub_wire78[719:704];
	wire [703:688] sub_wire76 = sub_wire1[703:688];
	wire [703:688] sub_wire75 = sub_wire76[703:688];
	wire [687:672] sub_wire74 = sub_wire1[687:672];
	wire [687:672] sub_wire73 = sub_wire74[687:672];
	wire [671:656] sub_wire72 = sub_wire1[671:656];
	wire [671:656] sub_wire71 = sub_wire72[671:656];
	wire [655:640] sub_wire70 = sub_wire1[655:640];
	wire [655:640] sub_wire69 = sub_wire70[655:640];
	wire [63:48] sub_wire68 = sub_wire1[63:48];
	wire [63:48] sub_wire67 = sub_wire68[63:48];
	wire [639:624] sub_wire66 = sub_wire1[639:624];
	wire [639:624] sub_wire65 = sub_wire66[639:624];
	wire [623:608] sub_wire64 = sub_wire1[623:608];
	wire [623:608] sub_wire63 = sub_wire64[623:608];
	wire [607:592] sub_wire62 = sub_wire1[607:592];
	wire [607:592] sub_wire61 = sub_wire62[607:592];
	wire [591:576] sub_wire60 = sub_wire1[591:576];
	wire [591:576] sub_wire59 = sub_wire60[591:576];
	wire [575:560] sub_wire58 = sub_wire1[575:560];
	wire [575:560] sub_wire57 = sub_wire58[575:560];
	wire [559:544] sub_wire56 = sub_wire1[559:544];
	wire [559:544] sub_wire55 = sub_wire56[559:544];
	wire [543:528] sub_wire54 = sub_wire1[543:528];
	wire [543:528] sub_wire53 = sub_wire54[543:528];
	wire [527:512] sub_wire52 = sub_wire1[527:512];
	wire [527:512] sub_wire51 = sub_wire52[527:512];
	wire [511:496] sub_wire50 = sub_wire1[511:496];
	wire [511:496] sub_wire49 = sub_wire50[511:496];
	wire [495:480] sub_wire48 = sub_wire1[495:480];
	wire [495:480] sub_wire47 = sub_wire48[495:480];
	wire [47:32] sub_wire46 = sub_wire1[47:32];
	wire [47:32] sub_wire45 = sub_wire46[47:32];
	wire [479:464] sub_wire44 = sub_wire1[479:464];
	wire [479:464] sub_wire43 = sub_wire44[479:464];
	wire [463:448] sub_wire42 = sub_wire1[463:448];
	wire [463:448] sub_wire41 = sub_wire42[463:448];
	wire [447:432] sub_wire40 = sub_wire1[447:432];
	wire [447:432] sub_wire39 = sub_wire40[447:432];
	wire [431:416] sub_wire38 = sub_wire1[431:416];
	wire [431:416] sub_wire37 = sub_wire38[431:416];
	wire [415:400] sub_wire36 = sub_wire1[415:400];
	wire [415:400] sub_wire35 = sub_wire36[415:400];
	wire [399:384] sub_wire34 = sub_wire1[399:384];
	wire [399:384] sub_wire33 = sub_wire34[399:384];
	wire [383:368] sub_wire32 = sub_wire1[383:368];
	wire [383:368] sub_wire31 = sub_wire32[383:368];
	wire [367:352] sub_wire30 = sub_wire1[367:352];
	wire [367:352] sub_wire29 = sub_wire30[367:352];
	wire [351:336] sub_wire28 = sub_wire1[351:336];
	wire [351:336] sub_wire27 = sub_wire28[351:336];
	wire [335:320] sub_wire26 = sub_wire1[335:320];
	wire [335:320] sub_wire25 = sub_wire26[335:320];
	wire [31:16] sub_wire24 = sub_wire1[31:16];
	wire [31:16] sub_wire23 = sub_wire24[31:16];
	wire [319:304] sub_wire22 = sub_wire1[319:304];
	wire [319:304] sub_wire21 = sub_wire22[319:304];
	wire [303:288] sub_wire20 = sub_wire1[303:288];
	wire [303:288] sub_wire19 = sub_wire20[303:288];
	wire [287:272] sub_wire18 = sub_wire1[287:272];
	wire [287:272] sub_wire17 = sub_wire18[287:272];
	wire [271:256] sub_wire16 = sub_wire1[271:256];
	wire [271:256] sub_wire15 = sub_wire16[271:256];
	wire [255:240] sub_wire14 = sub_wire1[255:240];
	wire [255:240] sub_wire13 = sub_wire14[255:240];
	wire [239:224] sub_wire12 = sub_wire1[239:224];
	wire [239:224] sub_wire11 = sub_wire12[239:224];
	wire [223:208] sub_wire10 = sub_wire1[223:208];
	wire [223:208] sub_wire9 = sub_wire10[223:208];
	wire [207:192] sub_wire8 = sub_wire1[207:192];
	wire [207:192] sub_wire7 = sub_wire8[207:192];
	wire [191:176] sub_wire6 = sub_wire1[191:176];
	wire [191:176] sub_wire5 = sub_wire6[191:176];
	wire [175:160] sub_wire4 = sub_wire1[175:160];
	wire [175:160] sub_wire3 = sub_wire4[175:160];
	wire [15:0] sub_wire2 = sub_wire1[15:0];
	wire [15:0] taps0x = sub_wire2[15:0];
	wire [15:0] taps10x = sub_wire3[175:160];
	wire [15:0] taps11x = sub_wire5[191:176];
	wire [15:0] taps12x = sub_wire7[207:192];
	wire [15:0] taps13x = sub_wire9[223:208];
	wire [15:0] taps14x = sub_wire11[239:224];
	wire [15:0] taps15x = sub_wire13[255:240];
	wire [15:0] taps16x = sub_wire15[271:256];
	wire [15:0] taps17x = sub_wire17[287:272];
	wire [15:0] taps18x = sub_wire19[303:288];
	wire [15:0] taps19x = sub_wire21[319:304];
	wire [15:0] taps1x = sub_wire23[31:16];
	wire [15:0] taps20x = sub_wire25[335:320];
	wire [15:0] taps21x = sub_wire27[351:336];
	wire [15:0] taps22x = sub_wire29[367:352];
	wire [15:0] taps23x = sub_wire31[383:368];
	wire [15:0] taps24x = sub_wire33[399:384];
	wire [15:0] taps25x = sub_wire35[415:400];
	wire [15:0] taps26x = sub_wire37[431:416];
	wire [15:0] taps27x = sub_wire39[447:432];
	wire [15:0] taps28x = sub_wire41[463:448];
	wire [15:0] taps29x = sub_wire43[479:464];
	wire [15:0] taps2x = sub_wire45[47:32];
	wire [15:0] taps30x = sub_wire47[495:480];
	wire [15:0] taps31x = sub_wire49[511:496];
	wire [15:0] taps32x = sub_wire51[527:512];
	wire [15:0] taps33x = sub_wire53[543:528];
	wire [15:0] taps34x = sub_wire55[559:544];
	wire [15:0] taps35x = sub_wire57[575:560];
	wire [15:0] taps36x = sub_wire59[591:576];
	wire [15:0] taps37x = sub_wire61[607:592];
	wire [15:0] taps38x = sub_wire63[623:608];
	wire [15:0] taps39x = sub_wire65[639:624];
	wire [15:0] taps3x = sub_wire67[63:48];
	wire [15:0] taps40x = sub_wire69[655:640];
	wire [15:0] taps41x = sub_wire71[671:656];
	wire [15:0] taps42x = sub_wire73[687:672];
	wire [15:0] taps43x = sub_wire75[703:688];
	wire [15:0] taps44x = sub_wire77[719:704];
	wire [15:0] taps45x = sub_wire79[735:720];
	wire [15:0] taps46x = sub_wire81[751:736];
	wire [15:0] taps47x = sub_wire83[767:752];
	wire [15:0] taps48x = sub_wire85[783:768];
	wire [15:0] taps49x = sub_wire87[799:784];
	wire [15:0] taps4x = sub_wire89[79:64];
	wire [15:0] taps50x = sub_wire91[815:800];
	wire [15:0] taps51x = sub_wire93[831:816];
	wire [15:0] taps52x = sub_wire95[847:832];
	wire [15:0] taps53x = sub_wire97[863:848];
	wire [15:0] taps54x = sub_wire99[879:864];
	wire [15:0] taps55x = sub_wire101[895:880];
	wire [15:0] taps56x = sub_wire103[911:896];
	wire [15:0] taps57x = sub_wire105[927:912];
	wire [15:0] taps58x = sub_wire107[943:928];
	wire [15:0] taps59x = sub_wire109[959:944];
	wire [15:0] taps5x = sub_wire111[95:80];
	wire [15:0] taps60x = sub_wire113[975:960];
	wire [15:0] taps61x = sub_wire115[991:976];
	wire [15:0] taps62x = sub_wire117[1007:992];
	wire [15:0] taps63x = sub_wire119[1023:1008];
	wire [15:0] taps64x = sub_wire121[1039:1024];
	wire [15:0] taps65x = sub_wire123[1055:1040];
	wire [15:0] taps66x = sub_wire125[1071:1056];
	wire [15:0] taps67x = sub_wire127[1087:1072];
	wire [15:0] taps68x = sub_wire129[1103:1088];
	wire [15:0] taps69x = sub_wire131[1119:1104];
	wire [15:0] taps6x = sub_wire133[111:96];
	wire [15:0] taps70x = sub_wire135[1135:1120];
	wire [15:0] taps71x = sub_wire137[1151:1136];
	wire [15:0] taps72x = sub_wire139[1167:1152];
	wire [15:0] taps73x = sub_wire141[1183:1168];
	wire [15:0] taps74x = sub_wire143[1199:1184];
	wire [15:0] taps75x = sub_wire145[1215:1200];
	wire [15:0] taps76x = sub_wire147[1231:1216];
	wire [15:0] taps77x = sub_wire149[1247:1232];
	wire [15:0] taps78x = sub_wire151[1263:1248];
	wire [15:0] taps79x = sub_wire153[1279:1264];
	wire [15:0] taps7x = sub_wire155[127:112];
	wire [15:0] taps80x = sub_wire157[1295:1280];
	wire [15:0] taps81x = sub_wire159[1311:1296];
	wire [15:0] taps82x = sub_wire161[1327:1312];
	wire [15:0] taps83x = sub_wire163[1343:1328];
	wire [15:0] taps84x = sub_wire165[1359:1344];
	wire [15:0] taps85x = sub_wire167[1375:1360];
	wire [15:0] taps86x = sub_wire169[1391:1376];
	wire [15:0] taps87x = sub_wire171[1407:1392];
	wire [15:0] taps88x = sub_wire173[1423:1408];
	wire [15:0] taps89x = sub_wire175[1439:1424];
	wire [15:0] taps8x = sub_wire177[143:128];
	wire [15:0] taps90x = sub_wire179[1455:1440];
	wire [15:0] taps91x = sub_wire181[1471:1456];
	wire [15:0] taps92x = sub_wire183[1487:1472];
	wire [15:0] taps93x = sub_wire185[1503:1488];
	wire [15:0] taps94x = sub_wire187[1519:1504];
	wire [15:0] taps95x = sub_wire189[1535:1520];
	wire [15:0] taps9x = sub_wire191[159:144];

	altshift_taps	ALTSHIFT_TAPS_component (
				.aclr (aclr),
				.clock (clock),
				.shiftin (shiftin),
				.shiftout (sub_wire0),
				.taps (sub_wire1)
				// synopsys translate_off
				,
				.clken (),
				.sclr ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Cyclone V",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 96,
		ALTSHIFT_TAPS_component.tap_distance = 4,
		ALTSHIFT_TAPS_component.width = 16;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "1"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "96"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "3"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "4"
// Retrieval info: PRIVATE: WIDTH NUMERIC "16"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=AUTO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "96"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "4"
// Retrieval info: CONSTANT: WIDTH NUMERIC "16"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT VCC "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 16 0 INPUT NODEFVAL "shiftin[15..0]"
// Retrieval info: USED_PORT: shiftout 0 0 16 0 OUTPUT NODEFVAL "shiftout[15..0]"
// Retrieval info: USED_PORT: taps0x 0 0 16 0 OUTPUT NODEFVAL "taps0x[15..0]"
// Retrieval info: USED_PORT: taps10x 0 0 16 0 OUTPUT NODEFVAL "taps10x[15..0]"
// Retrieval info: USED_PORT: taps11x 0 0 16 0 OUTPUT NODEFVAL "taps11x[15..0]"
// Retrieval info: USED_PORT: taps12x 0 0 16 0 OUTPUT NODEFVAL "taps12x[15..0]"
// Retrieval info: USED_PORT: taps13x 0 0 16 0 OUTPUT NODEFVAL "taps13x[15..0]"
// Retrieval info: USED_PORT: taps14x 0 0 16 0 OUTPUT NODEFVAL "taps14x[15..0]"
// Retrieval info: USED_PORT: taps15x 0 0 16 0 OUTPUT NODEFVAL "taps15x[15..0]"
// Retrieval info: USED_PORT: taps16x 0 0 16 0 OUTPUT NODEFVAL "taps16x[15..0]"
// Retrieval info: USED_PORT: taps17x 0 0 16 0 OUTPUT NODEFVAL "taps17x[15..0]"
// Retrieval info: USED_PORT: taps18x 0 0 16 0 OUTPUT NODEFVAL "taps18x[15..0]"
// Retrieval info: USED_PORT: taps19x 0 0 16 0 OUTPUT NODEFVAL "taps19x[15..0]"
// Retrieval info: USED_PORT: taps1x 0 0 16 0 OUTPUT NODEFVAL "taps1x[15..0]"
// Retrieval info: USED_PORT: taps20x 0 0 16 0 OUTPUT NODEFVAL "taps20x[15..0]"
// Retrieval info: USED_PORT: taps21x 0 0 16 0 OUTPUT NODEFVAL "taps21x[15..0]"
// Retrieval info: USED_PORT: taps22x 0 0 16 0 OUTPUT NODEFVAL "taps22x[15..0]"
// Retrieval info: USED_PORT: taps23x 0 0 16 0 OUTPUT NODEFVAL "taps23x[15..0]"
// Retrieval info: USED_PORT: taps24x 0 0 16 0 OUTPUT NODEFVAL "taps24x[15..0]"
// Retrieval info: USED_PORT: taps25x 0 0 16 0 OUTPUT NODEFVAL "taps25x[15..0]"
// Retrieval info: USED_PORT: taps26x 0 0 16 0 OUTPUT NODEFVAL "taps26x[15..0]"
// Retrieval info: USED_PORT: taps27x 0 0 16 0 OUTPUT NODEFVAL "taps27x[15..0]"
// Retrieval info: USED_PORT: taps28x 0 0 16 0 OUTPUT NODEFVAL "taps28x[15..0]"
// Retrieval info: USED_PORT: taps29x 0 0 16 0 OUTPUT NODEFVAL "taps29x[15..0]"
// Retrieval info: USED_PORT: taps2x 0 0 16 0 OUTPUT NODEFVAL "taps2x[15..0]"
// Retrieval info: USED_PORT: taps30x 0 0 16 0 OUTPUT NODEFVAL "taps30x[15..0]"
// Retrieval info: USED_PORT: taps31x 0 0 16 0 OUTPUT NODEFVAL "taps31x[15..0]"
// Retrieval info: USED_PORT: taps32x 0 0 16 0 OUTPUT NODEFVAL "taps32x[15..0]"
// Retrieval info: USED_PORT: taps33x 0 0 16 0 OUTPUT NODEFVAL "taps33x[15..0]"
// Retrieval info: USED_PORT: taps34x 0 0 16 0 OUTPUT NODEFVAL "taps34x[15..0]"
// Retrieval info: USED_PORT: taps35x 0 0 16 0 OUTPUT NODEFVAL "taps35x[15..0]"
// Retrieval info: USED_PORT: taps36x 0 0 16 0 OUTPUT NODEFVAL "taps36x[15..0]"
// Retrieval info: USED_PORT: taps37x 0 0 16 0 OUTPUT NODEFVAL "taps37x[15..0]"
// Retrieval info: USED_PORT: taps38x 0 0 16 0 OUTPUT NODEFVAL "taps38x[15..0]"
// Retrieval info: USED_PORT: taps39x 0 0 16 0 OUTPUT NODEFVAL "taps39x[15..0]"
// Retrieval info: USED_PORT: taps3x 0 0 16 0 OUTPUT NODEFVAL "taps3x[15..0]"
// Retrieval info: USED_PORT: taps40x 0 0 16 0 OUTPUT NODEFVAL "taps40x[15..0]"
// Retrieval info: USED_PORT: taps41x 0 0 16 0 OUTPUT NODEFVAL "taps41x[15..0]"
// Retrieval info: USED_PORT: taps42x 0 0 16 0 OUTPUT NODEFVAL "taps42x[15..0]"
// Retrieval info: USED_PORT: taps43x 0 0 16 0 OUTPUT NODEFVAL "taps43x[15..0]"
// Retrieval info: USED_PORT: taps44x 0 0 16 0 OUTPUT NODEFVAL "taps44x[15..0]"
// Retrieval info: USED_PORT: taps45x 0 0 16 0 OUTPUT NODEFVAL "taps45x[15..0]"
// Retrieval info: USED_PORT: taps46x 0 0 16 0 OUTPUT NODEFVAL "taps46x[15..0]"
// Retrieval info: USED_PORT: taps47x 0 0 16 0 OUTPUT NODEFVAL "taps47x[15..0]"
// Retrieval info: USED_PORT: taps48x 0 0 16 0 OUTPUT NODEFVAL "taps48x[15..0]"
// Retrieval info: USED_PORT: taps49x 0 0 16 0 OUTPUT NODEFVAL "taps49x[15..0]"
// Retrieval info: USED_PORT: taps4x 0 0 16 0 OUTPUT NODEFVAL "taps4x[15..0]"
// Retrieval info: USED_PORT: taps50x 0 0 16 0 OUTPUT NODEFVAL "taps50x[15..0]"
// Retrieval info: USED_PORT: taps51x 0 0 16 0 OUTPUT NODEFVAL "taps51x[15..0]"
// Retrieval info: USED_PORT: taps52x 0 0 16 0 OUTPUT NODEFVAL "taps52x[15..0]"
// Retrieval info: USED_PORT: taps53x 0 0 16 0 OUTPUT NODEFVAL "taps53x[15..0]"
// Retrieval info: USED_PORT: taps54x 0 0 16 0 OUTPUT NODEFVAL "taps54x[15..0]"
// Retrieval info: USED_PORT: taps55x 0 0 16 0 OUTPUT NODEFVAL "taps55x[15..0]"
// Retrieval info: USED_PORT: taps56x 0 0 16 0 OUTPUT NODEFVAL "taps56x[15..0]"
// Retrieval info: USED_PORT: taps57x 0 0 16 0 OUTPUT NODEFVAL "taps57x[15..0]"
// Retrieval info: USED_PORT: taps58x 0 0 16 0 OUTPUT NODEFVAL "taps58x[15..0]"
// Retrieval info: USED_PORT: taps59x 0 0 16 0 OUTPUT NODEFVAL "taps59x[15..0]"
// Retrieval info: USED_PORT: taps5x 0 0 16 0 OUTPUT NODEFVAL "taps5x[15..0]"
// Retrieval info: USED_PORT: taps60x 0 0 16 0 OUTPUT NODEFVAL "taps60x[15..0]"
// Retrieval info: USED_PORT: taps61x 0 0 16 0 OUTPUT NODEFVAL "taps61x[15..0]"
// Retrieval info: USED_PORT: taps62x 0 0 16 0 OUTPUT NODEFVAL "taps62x[15..0]"
// Retrieval info: USED_PORT: taps63x 0 0 16 0 OUTPUT NODEFVAL "taps63x[15..0]"
// Retrieval info: USED_PORT: taps64x 0 0 16 0 OUTPUT NODEFVAL "taps64x[15..0]"
// Retrieval info: USED_PORT: taps65x 0 0 16 0 OUTPUT NODEFVAL "taps65x[15..0]"
// Retrieval info: USED_PORT: taps66x 0 0 16 0 OUTPUT NODEFVAL "taps66x[15..0]"
// Retrieval info: USED_PORT: taps67x 0 0 16 0 OUTPUT NODEFVAL "taps67x[15..0]"
// Retrieval info: USED_PORT: taps68x 0 0 16 0 OUTPUT NODEFVAL "taps68x[15..0]"
// Retrieval info: USED_PORT: taps69x 0 0 16 0 OUTPUT NODEFVAL "taps69x[15..0]"
// Retrieval info: USED_PORT: taps6x 0 0 16 0 OUTPUT NODEFVAL "taps6x[15..0]"
// Retrieval info: USED_PORT: taps70x 0 0 16 0 OUTPUT NODEFVAL "taps70x[15..0]"
// Retrieval info: USED_PORT: taps71x 0 0 16 0 OUTPUT NODEFVAL "taps71x[15..0]"
// Retrieval info: USED_PORT: taps72x 0 0 16 0 OUTPUT NODEFVAL "taps72x[15..0]"
// Retrieval info: USED_PORT: taps73x 0 0 16 0 OUTPUT NODEFVAL "taps73x[15..0]"
// Retrieval info: USED_PORT: taps74x 0 0 16 0 OUTPUT NODEFVAL "taps74x[15..0]"
// Retrieval info: USED_PORT: taps75x 0 0 16 0 OUTPUT NODEFVAL "taps75x[15..0]"
// Retrieval info: USED_PORT: taps76x 0 0 16 0 OUTPUT NODEFVAL "taps76x[15..0]"
// Retrieval info: USED_PORT: taps77x 0 0 16 0 OUTPUT NODEFVAL "taps77x[15..0]"
// Retrieval info: USED_PORT: taps78x 0 0 16 0 OUTPUT NODEFVAL "taps78x[15..0]"
// Retrieval info: USED_PORT: taps79x 0 0 16 0 OUTPUT NODEFVAL "taps79x[15..0]"
// Retrieval info: USED_PORT: taps7x 0 0 16 0 OUTPUT NODEFVAL "taps7x[15..0]"
// Retrieval info: USED_PORT: taps80x 0 0 16 0 OUTPUT NODEFVAL "taps80x[15..0]"
// Retrieval info: USED_PORT: taps81x 0 0 16 0 OUTPUT NODEFVAL "taps81x[15..0]"
// Retrieval info: USED_PORT: taps82x 0 0 16 0 OUTPUT NODEFVAL "taps82x[15..0]"
// Retrieval info: USED_PORT: taps83x 0 0 16 0 OUTPUT NODEFVAL "taps83x[15..0]"
// Retrieval info: USED_PORT: taps84x 0 0 16 0 OUTPUT NODEFVAL "taps84x[15..0]"
// Retrieval info: USED_PORT: taps85x 0 0 16 0 OUTPUT NODEFVAL "taps85x[15..0]"
// Retrieval info: USED_PORT: taps86x 0 0 16 0 OUTPUT NODEFVAL "taps86x[15..0]"
// Retrieval info: USED_PORT: taps87x 0 0 16 0 OUTPUT NODEFVAL "taps87x[15..0]"
// Retrieval info: USED_PORT: taps88x 0 0 16 0 OUTPUT NODEFVAL "taps88x[15..0]"
// Retrieval info: USED_PORT: taps89x 0 0 16 0 OUTPUT NODEFVAL "taps89x[15..0]"
// Retrieval info: USED_PORT: taps8x 0 0 16 0 OUTPUT NODEFVAL "taps8x[15..0]"
// Retrieval info: USED_PORT: taps90x 0 0 16 0 OUTPUT NODEFVAL "taps90x[15..0]"
// Retrieval info: USED_PORT: taps91x 0 0 16 0 OUTPUT NODEFVAL "taps91x[15..0]"
// Retrieval info: USED_PORT: taps92x 0 0 16 0 OUTPUT NODEFVAL "taps92x[15..0]"
// Retrieval info: USED_PORT: taps93x 0 0 16 0 OUTPUT NODEFVAL "taps93x[15..0]"
// Retrieval info: USED_PORT: taps94x 0 0 16 0 OUTPUT NODEFVAL "taps94x[15..0]"
// Retrieval info: USED_PORT: taps95x 0 0 16 0 OUTPUT NODEFVAL "taps95x[15..0]"
// Retrieval info: USED_PORT: taps9x 0 0 16 0 OUTPUT NODEFVAL "taps9x[15..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 16 0 shiftin 0 0 16 0
// Retrieval info: CONNECT: shiftout 0 0 16 0 @shiftout 0 0 16 0
// Retrieval info: CONNECT: taps0x 0 0 16 0 @taps 0 0 16 0
// Retrieval info: CONNECT: taps10x 0 0 16 0 @taps 0 0 16 160
// Retrieval info: CONNECT: taps11x 0 0 16 0 @taps 0 0 16 176
// Retrieval info: CONNECT: taps12x 0 0 16 0 @taps 0 0 16 192
// Retrieval info: CONNECT: taps13x 0 0 16 0 @taps 0 0 16 208
// Retrieval info: CONNECT: taps14x 0 0 16 0 @taps 0 0 16 224
// Retrieval info: CONNECT: taps15x 0 0 16 0 @taps 0 0 16 240
// Retrieval info: CONNECT: taps16x 0 0 16 0 @taps 0 0 16 256
// Retrieval info: CONNECT: taps17x 0 0 16 0 @taps 0 0 16 272
// Retrieval info: CONNECT: taps18x 0 0 16 0 @taps 0 0 16 288
// Retrieval info: CONNECT: taps19x 0 0 16 0 @taps 0 0 16 304
// Retrieval info: CONNECT: taps1x 0 0 16 0 @taps 0 0 16 16
// Retrieval info: CONNECT: taps20x 0 0 16 0 @taps 0 0 16 320
// Retrieval info: CONNECT: taps21x 0 0 16 0 @taps 0 0 16 336
// Retrieval info: CONNECT: taps22x 0 0 16 0 @taps 0 0 16 352
// Retrieval info: CONNECT: taps23x 0 0 16 0 @taps 0 0 16 368
// Retrieval info: CONNECT: taps24x 0 0 16 0 @taps 0 0 16 384
// Retrieval info: CONNECT: taps25x 0 0 16 0 @taps 0 0 16 400
// Retrieval info: CONNECT: taps26x 0 0 16 0 @taps 0 0 16 416
// Retrieval info: CONNECT: taps27x 0 0 16 0 @taps 0 0 16 432
// Retrieval info: CONNECT: taps28x 0 0 16 0 @taps 0 0 16 448
// Retrieval info: CONNECT: taps29x 0 0 16 0 @taps 0 0 16 464
// Retrieval info: CONNECT: taps2x 0 0 16 0 @taps 0 0 16 32
// Retrieval info: CONNECT: taps30x 0 0 16 0 @taps 0 0 16 480
// Retrieval info: CONNECT: taps31x 0 0 16 0 @taps 0 0 16 496
// Retrieval info: CONNECT: taps32x 0 0 16 0 @taps 0 0 16 512
// Retrieval info: CONNECT: taps33x 0 0 16 0 @taps 0 0 16 528
// Retrieval info: CONNECT: taps34x 0 0 16 0 @taps 0 0 16 544
// Retrieval info: CONNECT: taps35x 0 0 16 0 @taps 0 0 16 560
// Retrieval info: CONNECT: taps36x 0 0 16 0 @taps 0 0 16 576
// Retrieval info: CONNECT: taps37x 0 0 16 0 @taps 0 0 16 592
// Retrieval info: CONNECT: taps38x 0 0 16 0 @taps 0 0 16 608
// Retrieval info: CONNECT: taps39x 0 0 16 0 @taps 0 0 16 624
// Retrieval info: CONNECT: taps3x 0 0 16 0 @taps 0 0 16 48
// Retrieval info: CONNECT: taps40x 0 0 16 0 @taps 0 0 16 640
// Retrieval info: CONNECT: taps41x 0 0 16 0 @taps 0 0 16 656
// Retrieval info: CONNECT: taps42x 0 0 16 0 @taps 0 0 16 672
// Retrieval info: CONNECT: taps43x 0 0 16 0 @taps 0 0 16 688
// Retrieval info: CONNECT: taps44x 0 0 16 0 @taps 0 0 16 704
// Retrieval info: CONNECT: taps45x 0 0 16 0 @taps 0 0 16 720
// Retrieval info: CONNECT: taps46x 0 0 16 0 @taps 0 0 16 736
// Retrieval info: CONNECT: taps47x 0 0 16 0 @taps 0 0 16 752
// Retrieval info: CONNECT: taps48x 0 0 16 0 @taps 0 0 16 768
// Retrieval info: CONNECT: taps49x 0 0 16 0 @taps 0 0 16 784
// Retrieval info: CONNECT: taps4x 0 0 16 0 @taps 0 0 16 64
// Retrieval info: CONNECT: taps50x 0 0 16 0 @taps 0 0 16 800
// Retrieval info: CONNECT: taps51x 0 0 16 0 @taps 0 0 16 816
// Retrieval info: CONNECT: taps52x 0 0 16 0 @taps 0 0 16 832
// Retrieval info: CONNECT: taps53x 0 0 16 0 @taps 0 0 16 848
// Retrieval info: CONNECT: taps54x 0 0 16 0 @taps 0 0 16 864
// Retrieval info: CONNECT: taps55x 0 0 16 0 @taps 0 0 16 880
// Retrieval info: CONNECT: taps56x 0 0 16 0 @taps 0 0 16 896
// Retrieval info: CONNECT: taps57x 0 0 16 0 @taps 0 0 16 912
// Retrieval info: CONNECT: taps58x 0 0 16 0 @taps 0 0 16 928
// Retrieval info: CONNECT: taps59x 0 0 16 0 @taps 0 0 16 944
// Retrieval info: CONNECT: taps5x 0 0 16 0 @taps 0 0 16 80
// Retrieval info: CONNECT: taps60x 0 0 16 0 @taps 0 0 16 960
// Retrieval info: CONNECT: taps61x 0 0 16 0 @taps 0 0 16 976
// Retrieval info: CONNECT: taps62x 0 0 16 0 @taps 0 0 16 992
// Retrieval info: CONNECT: taps63x 0 0 16 0 @taps 0 0 16 1008
// Retrieval info: CONNECT: taps64x 0 0 16 0 @taps 0 0 16 1024
// Retrieval info: CONNECT: taps65x 0 0 16 0 @taps 0 0 16 1040
// Retrieval info: CONNECT: taps66x 0 0 16 0 @taps 0 0 16 1056
// Retrieval info: CONNECT: taps67x 0 0 16 0 @taps 0 0 16 1072
// Retrieval info: CONNECT: taps68x 0 0 16 0 @taps 0 0 16 1088
// Retrieval info: CONNECT: taps69x 0 0 16 0 @taps 0 0 16 1104
// Retrieval info: CONNECT: taps6x 0 0 16 0 @taps 0 0 16 96
// Retrieval info: CONNECT: taps70x 0 0 16 0 @taps 0 0 16 1120
// Retrieval info: CONNECT: taps71x 0 0 16 0 @taps 0 0 16 1136
// Retrieval info: CONNECT: taps72x 0 0 16 0 @taps 0 0 16 1152
// Retrieval info: CONNECT: taps73x 0 0 16 0 @taps 0 0 16 1168
// Retrieval info: CONNECT: taps74x 0 0 16 0 @taps 0 0 16 1184
// Retrieval info: CONNECT: taps75x 0 0 16 0 @taps 0 0 16 1200
// Retrieval info: CONNECT: taps76x 0 0 16 0 @taps 0 0 16 1216
// Retrieval info: CONNECT: taps77x 0 0 16 0 @taps 0 0 16 1232
// Retrieval info: CONNECT: taps78x 0 0 16 0 @taps 0 0 16 1248
// Retrieval info: CONNECT: taps79x 0 0 16 0 @taps 0 0 16 1264
// Retrieval info: CONNECT: taps7x 0 0 16 0 @taps 0 0 16 112
// Retrieval info: CONNECT: taps80x 0 0 16 0 @taps 0 0 16 1280
// Retrieval info: CONNECT: taps81x 0 0 16 0 @taps 0 0 16 1296
// Retrieval info: CONNECT: taps82x 0 0 16 0 @taps 0 0 16 1312
// Retrieval info: CONNECT: taps83x 0 0 16 0 @taps 0 0 16 1328
// Retrieval info: CONNECT: taps84x 0 0 16 0 @taps 0 0 16 1344
// Retrieval info: CONNECT: taps85x 0 0 16 0 @taps 0 0 16 1360
// Retrieval info: CONNECT: taps86x 0 0 16 0 @taps 0 0 16 1376
// Retrieval info: CONNECT: taps87x 0 0 16 0 @taps 0 0 16 1392
// Retrieval info: CONNECT: taps88x 0 0 16 0 @taps 0 0 16 1408
// Retrieval info: CONNECT: taps89x 0 0 16 0 @taps 0 0 16 1424
// Retrieval info: CONNECT: taps8x 0 0 16 0 @taps 0 0 16 128
// Retrieval info: CONNECT: taps90x 0 0 16 0 @taps 0 0 16 1440
// Retrieval info: CONNECT: taps91x 0 0 16 0 @taps 0 0 16 1456
// Retrieval info: CONNECT: taps92x 0 0 16 0 @taps 0 0 16 1472
// Retrieval info: CONNECT: taps93x 0 0 16 0 @taps 0 0 16 1488
// Retrieval info: CONNECT: taps94x 0 0 16 0 @taps 0 0 16 1504
// Retrieval info: CONNECT: taps95x 0 0 16 0 @taps 0 0 16 1520
// Retrieval info: CONNECT: taps9x 0 0 16 0 @taps 0 0 16 144
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
