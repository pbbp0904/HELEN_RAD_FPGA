// megafunction wizard: %Shift register (RAM-based)%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: Shift.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************

//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module Shift (
	aclr,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps10x,
	taps11x,
	taps12x,
	taps13x,
	taps14x,
	taps15x,
	taps16x,
	taps17x,
	taps18x,
	taps19x,
	taps1x,
	taps20x,
	taps21x,
	taps22x,
	taps23x,
	taps24x,
	taps25x,
	taps26x,
	taps27x,
	taps28x,
	taps29x,
	taps2x,
	taps30x,
	taps31x,
	taps32x,
	taps33x,
	taps34x,
	taps35x,
	taps36x,
	taps37x,
	taps38x,
	taps39x,
	taps3x,
	taps40x,
	taps41x,
	taps42x,
	taps43x,
	taps44x,
	taps45x,
	taps46x,
	taps47x,
	taps48x,
	taps49x,
	taps4x,
	taps50x,
	taps51x,
	taps52x,
	taps53x,
	taps54x,
	taps55x,
	taps56x,
	taps57x,
	taps58x,
	taps59x,
	taps5x,
	taps60x,
	taps61x,
	taps62x,
	taps63x,
	taps64x,
	taps65x,
	taps66x,
	taps67x,
	taps68x,
	taps69x,
	taps6x,
	taps70x,
	taps71x,
	taps72x,
	taps73x,
	taps74x,
	taps75x,
	taps76x,
	taps77x,
	taps78x,
	taps79x,
	taps7x,
	taps80x,
	taps81x,
	taps82x,
	taps83x,
	taps84x,
	taps85x,
	taps86x,
	taps87x,
	taps88x,
	taps89x,
	taps8x,
	taps90x,
	taps91x,
	taps92x,
	taps93x,
	taps94x,
	taps95x,
	taps9x);

	input	  aclr;
	input	  clock;
	input	[15:0]  shiftin;
	output	[15:0]  shiftout;
	output	[15:0]  taps0x;
	output	[15:0]  taps10x;
	output	[15:0]  taps11x;
	output	[15:0]  taps12x;
	output	[15:0]  taps13x;
	output	[15:0]  taps14x;
	output	[15:0]  taps15x;
	output	[15:0]  taps16x;
	output	[15:0]  taps17x;
	output	[15:0]  taps18x;
	output	[15:0]  taps19x;
	output	[15:0]  taps1x;
	output	[15:0]  taps20x;
	output	[15:0]  taps21x;
	output	[15:0]  taps22x;
	output	[15:0]  taps23x;
	output	[15:0]  taps24x;
	output	[15:0]  taps25x;
	output	[15:0]  taps26x;
	output	[15:0]  taps27x;
	output	[15:0]  taps28x;
	output	[15:0]  taps29x;
	output	[15:0]  taps2x;
	output	[15:0]  taps30x;
	output	[15:0]  taps31x;
	output	[15:0]  taps32x;
	output	[15:0]  taps33x;
	output	[15:0]  taps34x;
	output	[15:0]  taps35x;
	output	[15:0]  taps36x;
	output	[15:0]  taps37x;
	output	[15:0]  taps38x;
	output	[15:0]  taps39x;
	output	[15:0]  taps3x;
	output	[15:0]  taps40x;
	output	[15:0]  taps41x;
	output	[15:0]  taps42x;
	output	[15:0]  taps43x;
	output	[15:0]  taps44x;
	output	[15:0]  taps45x;
	output	[15:0]  taps46x;
	output	[15:0]  taps47x;
	output	[15:0]  taps48x;
	output	[15:0]  taps49x;
	output	[15:0]  taps4x;
	output	[15:0]  taps50x;
	output	[15:0]  taps51x;
	output	[15:0]  taps52x;
	output	[15:0]  taps53x;
	output	[15:0]  taps54x;
	output	[15:0]  taps55x;
	output	[15:0]  taps56x;
	output	[15:0]  taps57x;
	output	[15:0]  taps58x;
	output	[15:0]  taps59x;
	output	[15:0]  taps5x;
	output	[15:0]  taps60x;
	output	[15:0]  taps61x;
	output	[15:0]  taps62x;
	output	[15:0]  taps63x;
	output	[15:0]  taps64x;
	output	[15:0]  taps65x;
	output	[15:0]  taps66x;
	output	[15:0]  taps67x;
	output	[15:0]  taps68x;
	output	[15:0]  taps69x;
	output	[15:0]  taps6x;
	output	[15:0]  taps70x;
	output	[15:0]  taps71x;
	output	[15:0]  taps72x;
	output	[15:0]  taps73x;
	output	[15:0]  taps74x;
	output	[15:0]  taps75x;
	output	[15:0]  taps76x;
	output	[15:0]  taps77x;
	output	[15:0]  taps78x;
	output	[15:0]  taps79x;
	output	[15:0]  taps7x;
	output	[15:0]  taps80x;
	output	[15:0]  taps81x;
	output	[15:0]  taps82x;
	output	[15:0]  taps83x;
	output	[15:0]  taps84x;
	output	[15:0]  taps85x;
	output	[15:0]  taps86x;
	output	[15:0]  taps87x;
	output	[15:0]  taps88x;
	output	[15:0]  taps89x;
	output	[15:0]  taps8x;
	output	[15:0]  taps90x;
	output	[15:0]  taps91x;
	output	[15:0]  taps92x;
	output	[15:0]  taps93x;
	output	[15:0]  taps94x;
	output	[15:0]  taps95x;
	output	[15:0]  taps9x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  aclr;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "1"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "96"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "3"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "4"
// Retrieval info: PRIVATE: WIDTH NUMERIC "16"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=AUTO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "96"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "4"
// Retrieval info: CONSTANT: WIDTH NUMERIC "16"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT VCC "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 16 0 INPUT NODEFVAL "shiftin[15..0]"
// Retrieval info: USED_PORT: shiftout 0 0 16 0 OUTPUT NODEFVAL "shiftout[15..0]"
// Retrieval info: USED_PORT: taps0x 0 0 16 0 OUTPUT NODEFVAL "taps0x[15..0]"
// Retrieval info: USED_PORT: taps10x 0 0 16 0 OUTPUT NODEFVAL "taps10x[15..0]"
// Retrieval info: USED_PORT: taps11x 0 0 16 0 OUTPUT NODEFVAL "taps11x[15..0]"
// Retrieval info: USED_PORT: taps12x 0 0 16 0 OUTPUT NODEFVAL "taps12x[15..0]"
// Retrieval info: USED_PORT: taps13x 0 0 16 0 OUTPUT NODEFVAL "taps13x[15..0]"
// Retrieval info: USED_PORT: taps14x 0 0 16 0 OUTPUT NODEFVAL "taps14x[15..0]"
// Retrieval info: USED_PORT: taps15x 0 0 16 0 OUTPUT NODEFVAL "taps15x[15..0]"
// Retrieval info: USED_PORT: taps16x 0 0 16 0 OUTPUT NODEFVAL "taps16x[15..0]"
// Retrieval info: USED_PORT: taps17x 0 0 16 0 OUTPUT NODEFVAL "taps17x[15..0]"
// Retrieval info: USED_PORT: taps18x 0 0 16 0 OUTPUT NODEFVAL "taps18x[15..0]"
// Retrieval info: USED_PORT: taps19x 0 0 16 0 OUTPUT NODEFVAL "taps19x[15..0]"
// Retrieval info: USED_PORT: taps1x 0 0 16 0 OUTPUT NODEFVAL "taps1x[15..0]"
// Retrieval info: USED_PORT: taps20x 0 0 16 0 OUTPUT NODEFVAL "taps20x[15..0]"
// Retrieval info: USED_PORT: taps21x 0 0 16 0 OUTPUT NODEFVAL "taps21x[15..0]"
// Retrieval info: USED_PORT: taps22x 0 0 16 0 OUTPUT NODEFVAL "taps22x[15..0]"
// Retrieval info: USED_PORT: taps23x 0 0 16 0 OUTPUT NODEFVAL "taps23x[15..0]"
// Retrieval info: USED_PORT: taps24x 0 0 16 0 OUTPUT NODEFVAL "taps24x[15..0]"
// Retrieval info: USED_PORT: taps25x 0 0 16 0 OUTPUT NODEFVAL "taps25x[15..0]"
// Retrieval info: USED_PORT: taps26x 0 0 16 0 OUTPUT NODEFVAL "taps26x[15..0]"
// Retrieval info: USED_PORT: taps27x 0 0 16 0 OUTPUT NODEFVAL "taps27x[15..0]"
// Retrieval info: USED_PORT: taps28x 0 0 16 0 OUTPUT NODEFVAL "taps28x[15..0]"
// Retrieval info: USED_PORT: taps29x 0 0 16 0 OUTPUT NODEFVAL "taps29x[15..0]"
// Retrieval info: USED_PORT: taps2x 0 0 16 0 OUTPUT NODEFVAL "taps2x[15..0]"
// Retrieval info: USED_PORT: taps30x 0 0 16 0 OUTPUT NODEFVAL "taps30x[15..0]"
// Retrieval info: USED_PORT: taps31x 0 0 16 0 OUTPUT NODEFVAL "taps31x[15..0]"
// Retrieval info: USED_PORT: taps32x 0 0 16 0 OUTPUT NODEFVAL "taps32x[15..0]"
// Retrieval info: USED_PORT: taps33x 0 0 16 0 OUTPUT NODEFVAL "taps33x[15..0]"
// Retrieval info: USED_PORT: taps34x 0 0 16 0 OUTPUT NODEFVAL "taps34x[15..0]"
// Retrieval info: USED_PORT: taps35x 0 0 16 0 OUTPUT NODEFVAL "taps35x[15..0]"
// Retrieval info: USED_PORT: taps36x 0 0 16 0 OUTPUT NODEFVAL "taps36x[15..0]"
// Retrieval info: USED_PORT: taps37x 0 0 16 0 OUTPUT NODEFVAL "taps37x[15..0]"
// Retrieval info: USED_PORT: taps38x 0 0 16 0 OUTPUT NODEFVAL "taps38x[15..0]"
// Retrieval info: USED_PORT: taps39x 0 0 16 0 OUTPUT NODEFVAL "taps39x[15..0]"
// Retrieval info: USED_PORT: taps3x 0 0 16 0 OUTPUT NODEFVAL "taps3x[15..0]"
// Retrieval info: USED_PORT: taps40x 0 0 16 0 OUTPUT NODEFVAL "taps40x[15..0]"
// Retrieval info: USED_PORT: taps41x 0 0 16 0 OUTPUT NODEFVAL "taps41x[15..0]"
// Retrieval info: USED_PORT: taps42x 0 0 16 0 OUTPUT NODEFVAL "taps42x[15..0]"
// Retrieval info: USED_PORT: taps43x 0 0 16 0 OUTPUT NODEFVAL "taps43x[15..0]"
// Retrieval info: USED_PORT: taps44x 0 0 16 0 OUTPUT NODEFVAL "taps44x[15..0]"
// Retrieval info: USED_PORT: taps45x 0 0 16 0 OUTPUT NODEFVAL "taps45x[15..0]"
// Retrieval info: USED_PORT: taps46x 0 0 16 0 OUTPUT NODEFVAL "taps46x[15..0]"
// Retrieval info: USED_PORT: taps47x 0 0 16 0 OUTPUT NODEFVAL "taps47x[15..0]"
// Retrieval info: USED_PORT: taps48x 0 0 16 0 OUTPUT NODEFVAL "taps48x[15..0]"
// Retrieval info: USED_PORT: taps49x 0 0 16 0 OUTPUT NODEFVAL "taps49x[15..0]"
// Retrieval info: USED_PORT: taps4x 0 0 16 0 OUTPUT NODEFVAL "taps4x[15..0]"
// Retrieval info: USED_PORT: taps50x 0 0 16 0 OUTPUT NODEFVAL "taps50x[15..0]"
// Retrieval info: USED_PORT: taps51x 0 0 16 0 OUTPUT NODEFVAL "taps51x[15..0]"
// Retrieval info: USED_PORT: taps52x 0 0 16 0 OUTPUT NODEFVAL "taps52x[15..0]"
// Retrieval info: USED_PORT: taps53x 0 0 16 0 OUTPUT NODEFVAL "taps53x[15..0]"
// Retrieval info: USED_PORT: taps54x 0 0 16 0 OUTPUT NODEFVAL "taps54x[15..0]"
// Retrieval info: USED_PORT: taps55x 0 0 16 0 OUTPUT NODEFVAL "taps55x[15..0]"
// Retrieval info: USED_PORT: taps56x 0 0 16 0 OUTPUT NODEFVAL "taps56x[15..0]"
// Retrieval info: USED_PORT: taps57x 0 0 16 0 OUTPUT NODEFVAL "taps57x[15..0]"
// Retrieval info: USED_PORT: taps58x 0 0 16 0 OUTPUT NODEFVAL "taps58x[15..0]"
// Retrieval info: USED_PORT: taps59x 0 0 16 0 OUTPUT NODEFVAL "taps59x[15..0]"
// Retrieval info: USED_PORT: taps5x 0 0 16 0 OUTPUT NODEFVAL "taps5x[15..0]"
// Retrieval info: USED_PORT: taps60x 0 0 16 0 OUTPUT NODEFVAL "taps60x[15..0]"
// Retrieval info: USED_PORT: taps61x 0 0 16 0 OUTPUT NODEFVAL "taps61x[15..0]"
// Retrieval info: USED_PORT: taps62x 0 0 16 0 OUTPUT NODEFVAL "taps62x[15..0]"
// Retrieval info: USED_PORT: taps63x 0 0 16 0 OUTPUT NODEFVAL "taps63x[15..0]"
// Retrieval info: USED_PORT: taps64x 0 0 16 0 OUTPUT NODEFVAL "taps64x[15..0]"
// Retrieval info: USED_PORT: taps65x 0 0 16 0 OUTPUT NODEFVAL "taps65x[15..0]"
// Retrieval info: USED_PORT: taps66x 0 0 16 0 OUTPUT NODEFVAL "taps66x[15..0]"
// Retrieval info: USED_PORT: taps67x 0 0 16 0 OUTPUT NODEFVAL "taps67x[15..0]"
// Retrieval info: USED_PORT: taps68x 0 0 16 0 OUTPUT NODEFVAL "taps68x[15..0]"
// Retrieval info: USED_PORT: taps69x 0 0 16 0 OUTPUT NODEFVAL "taps69x[15..0]"
// Retrieval info: USED_PORT: taps6x 0 0 16 0 OUTPUT NODEFVAL "taps6x[15..0]"
// Retrieval info: USED_PORT: taps70x 0 0 16 0 OUTPUT NODEFVAL "taps70x[15..0]"
// Retrieval info: USED_PORT: taps71x 0 0 16 0 OUTPUT NODEFVAL "taps71x[15..0]"
// Retrieval info: USED_PORT: taps72x 0 0 16 0 OUTPUT NODEFVAL "taps72x[15..0]"
// Retrieval info: USED_PORT: taps73x 0 0 16 0 OUTPUT NODEFVAL "taps73x[15..0]"
// Retrieval info: USED_PORT: taps74x 0 0 16 0 OUTPUT NODEFVAL "taps74x[15..0]"
// Retrieval info: USED_PORT: taps75x 0 0 16 0 OUTPUT NODEFVAL "taps75x[15..0]"
// Retrieval info: USED_PORT: taps76x 0 0 16 0 OUTPUT NODEFVAL "taps76x[15..0]"
// Retrieval info: USED_PORT: taps77x 0 0 16 0 OUTPUT NODEFVAL "taps77x[15..0]"
// Retrieval info: USED_PORT: taps78x 0 0 16 0 OUTPUT NODEFVAL "taps78x[15..0]"
// Retrieval info: USED_PORT: taps79x 0 0 16 0 OUTPUT NODEFVAL "taps79x[15..0]"
// Retrieval info: USED_PORT: taps7x 0 0 16 0 OUTPUT NODEFVAL "taps7x[15..0]"
// Retrieval info: USED_PORT: taps80x 0 0 16 0 OUTPUT NODEFVAL "taps80x[15..0]"
// Retrieval info: USED_PORT: taps81x 0 0 16 0 OUTPUT NODEFVAL "taps81x[15..0]"
// Retrieval info: USED_PORT: taps82x 0 0 16 0 OUTPUT NODEFVAL "taps82x[15..0]"
// Retrieval info: USED_PORT: taps83x 0 0 16 0 OUTPUT NODEFVAL "taps83x[15..0]"
// Retrieval info: USED_PORT: taps84x 0 0 16 0 OUTPUT NODEFVAL "taps84x[15..0]"
// Retrieval info: USED_PORT: taps85x 0 0 16 0 OUTPUT NODEFVAL "taps85x[15..0]"
// Retrieval info: USED_PORT: taps86x 0 0 16 0 OUTPUT NODEFVAL "taps86x[15..0]"
// Retrieval info: USED_PORT: taps87x 0 0 16 0 OUTPUT NODEFVAL "taps87x[15..0]"
// Retrieval info: USED_PORT: taps88x 0 0 16 0 OUTPUT NODEFVAL "taps88x[15..0]"
// Retrieval info: USED_PORT: taps89x 0 0 16 0 OUTPUT NODEFVAL "taps89x[15..0]"
// Retrieval info: USED_PORT: taps8x 0 0 16 0 OUTPUT NODEFVAL "taps8x[15..0]"
// Retrieval info: USED_PORT: taps90x 0 0 16 0 OUTPUT NODEFVAL "taps90x[15..0]"
// Retrieval info: USED_PORT: taps91x 0 0 16 0 OUTPUT NODEFVAL "taps91x[15..0]"
// Retrieval info: USED_PORT: taps92x 0 0 16 0 OUTPUT NODEFVAL "taps92x[15..0]"
// Retrieval info: USED_PORT: taps93x 0 0 16 0 OUTPUT NODEFVAL "taps93x[15..0]"
// Retrieval info: USED_PORT: taps94x 0 0 16 0 OUTPUT NODEFVAL "taps94x[15..0]"
// Retrieval info: USED_PORT: taps95x 0 0 16 0 OUTPUT NODEFVAL "taps95x[15..0]"
// Retrieval info: USED_PORT: taps9x 0 0 16 0 OUTPUT NODEFVAL "taps9x[15..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 16 0 shiftin 0 0 16 0
// Retrieval info: CONNECT: shiftout 0 0 16 0 @shiftout 0 0 16 0
// Retrieval info: CONNECT: taps0x 0 0 16 0 @taps 0 0 16 0
// Retrieval info: CONNECT: taps10x 0 0 16 0 @taps 0 0 16 160
// Retrieval info: CONNECT: taps11x 0 0 16 0 @taps 0 0 16 176
// Retrieval info: CONNECT: taps12x 0 0 16 0 @taps 0 0 16 192
// Retrieval info: CONNECT: taps13x 0 0 16 0 @taps 0 0 16 208
// Retrieval info: CONNECT: taps14x 0 0 16 0 @taps 0 0 16 224
// Retrieval info: CONNECT: taps15x 0 0 16 0 @taps 0 0 16 240
// Retrieval info: CONNECT: taps16x 0 0 16 0 @taps 0 0 16 256
// Retrieval info: CONNECT: taps17x 0 0 16 0 @taps 0 0 16 272
// Retrieval info: CONNECT: taps18x 0 0 16 0 @taps 0 0 16 288
// Retrieval info: CONNECT: taps19x 0 0 16 0 @taps 0 0 16 304
// Retrieval info: CONNECT: taps1x 0 0 16 0 @taps 0 0 16 16
// Retrieval info: CONNECT: taps20x 0 0 16 0 @taps 0 0 16 320
// Retrieval info: CONNECT: taps21x 0 0 16 0 @taps 0 0 16 336
// Retrieval info: CONNECT: taps22x 0 0 16 0 @taps 0 0 16 352
// Retrieval info: CONNECT: taps23x 0 0 16 0 @taps 0 0 16 368
// Retrieval info: CONNECT: taps24x 0 0 16 0 @taps 0 0 16 384
// Retrieval info: CONNECT: taps25x 0 0 16 0 @taps 0 0 16 400
// Retrieval info: CONNECT: taps26x 0 0 16 0 @taps 0 0 16 416
// Retrieval info: CONNECT: taps27x 0 0 16 0 @taps 0 0 16 432
// Retrieval info: CONNECT: taps28x 0 0 16 0 @taps 0 0 16 448
// Retrieval info: CONNECT: taps29x 0 0 16 0 @taps 0 0 16 464
// Retrieval info: CONNECT: taps2x 0 0 16 0 @taps 0 0 16 32
// Retrieval info: CONNECT: taps30x 0 0 16 0 @taps 0 0 16 480
// Retrieval info: CONNECT: taps31x 0 0 16 0 @taps 0 0 16 496
// Retrieval info: CONNECT: taps32x 0 0 16 0 @taps 0 0 16 512
// Retrieval info: CONNECT: taps33x 0 0 16 0 @taps 0 0 16 528
// Retrieval info: CONNECT: taps34x 0 0 16 0 @taps 0 0 16 544
// Retrieval info: CONNECT: taps35x 0 0 16 0 @taps 0 0 16 560
// Retrieval info: CONNECT: taps36x 0 0 16 0 @taps 0 0 16 576
// Retrieval info: CONNECT: taps37x 0 0 16 0 @taps 0 0 16 592
// Retrieval info: CONNECT: taps38x 0 0 16 0 @taps 0 0 16 608
// Retrieval info: CONNECT: taps39x 0 0 16 0 @taps 0 0 16 624
// Retrieval info: CONNECT: taps3x 0 0 16 0 @taps 0 0 16 48
// Retrieval info: CONNECT: taps40x 0 0 16 0 @taps 0 0 16 640
// Retrieval info: CONNECT: taps41x 0 0 16 0 @taps 0 0 16 656
// Retrieval info: CONNECT: taps42x 0 0 16 0 @taps 0 0 16 672
// Retrieval info: CONNECT: taps43x 0 0 16 0 @taps 0 0 16 688
// Retrieval info: CONNECT: taps44x 0 0 16 0 @taps 0 0 16 704
// Retrieval info: CONNECT: taps45x 0 0 16 0 @taps 0 0 16 720
// Retrieval info: CONNECT: taps46x 0 0 16 0 @taps 0 0 16 736
// Retrieval info: CONNECT: taps47x 0 0 16 0 @taps 0 0 16 752
// Retrieval info: CONNECT: taps48x 0 0 16 0 @taps 0 0 16 768
// Retrieval info: CONNECT: taps49x 0 0 16 0 @taps 0 0 16 784
// Retrieval info: CONNECT: taps4x 0 0 16 0 @taps 0 0 16 64
// Retrieval info: CONNECT: taps50x 0 0 16 0 @taps 0 0 16 800
// Retrieval info: CONNECT: taps51x 0 0 16 0 @taps 0 0 16 816
// Retrieval info: CONNECT: taps52x 0 0 16 0 @taps 0 0 16 832
// Retrieval info: CONNECT: taps53x 0 0 16 0 @taps 0 0 16 848
// Retrieval info: CONNECT: taps54x 0 0 16 0 @taps 0 0 16 864
// Retrieval info: CONNECT: taps55x 0 0 16 0 @taps 0 0 16 880
// Retrieval info: CONNECT: taps56x 0 0 16 0 @taps 0 0 16 896
// Retrieval info: CONNECT: taps57x 0 0 16 0 @taps 0 0 16 912
// Retrieval info: CONNECT: taps58x 0 0 16 0 @taps 0 0 16 928
// Retrieval info: CONNECT: taps59x 0 0 16 0 @taps 0 0 16 944
// Retrieval info: CONNECT: taps5x 0 0 16 0 @taps 0 0 16 80
// Retrieval info: CONNECT: taps60x 0 0 16 0 @taps 0 0 16 960
// Retrieval info: CONNECT: taps61x 0 0 16 0 @taps 0 0 16 976
// Retrieval info: CONNECT: taps62x 0 0 16 0 @taps 0 0 16 992
// Retrieval info: CONNECT: taps63x 0 0 16 0 @taps 0 0 16 1008
// Retrieval info: CONNECT: taps64x 0 0 16 0 @taps 0 0 16 1024
// Retrieval info: CONNECT: taps65x 0 0 16 0 @taps 0 0 16 1040
// Retrieval info: CONNECT: taps66x 0 0 16 0 @taps 0 0 16 1056
// Retrieval info: CONNECT: taps67x 0 0 16 0 @taps 0 0 16 1072
// Retrieval info: CONNECT: taps68x 0 0 16 0 @taps 0 0 16 1088
// Retrieval info: CONNECT: taps69x 0 0 16 0 @taps 0 0 16 1104
// Retrieval info: CONNECT: taps6x 0 0 16 0 @taps 0 0 16 96
// Retrieval info: CONNECT: taps70x 0 0 16 0 @taps 0 0 16 1120
// Retrieval info: CONNECT: taps71x 0 0 16 0 @taps 0 0 16 1136
// Retrieval info: CONNECT: taps72x 0 0 16 0 @taps 0 0 16 1152
// Retrieval info: CONNECT: taps73x 0 0 16 0 @taps 0 0 16 1168
// Retrieval info: CONNECT: taps74x 0 0 16 0 @taps 0 0 16 1184
// Retrieval info: CONNECT: taps75x 0 0 16 0 @taps 0 0 16 1200
// Retrieval info: CONNECT: taps76x 0 0 16 0 @taps 0 0 16 1216
// Retrieval info: CONNECT: taps77x 0 0 16 0 @taps 0 0 16 1232
// Retrieval info: CONNECT: taps78x 0 0 16 0 @taps 0 0 16 1248
// Retrieval info: CONNECT: taps79x 0 0 16 0 @taps 0 0 16 1264
// Retrieval info: CONNECT: taps7x 0 0 16 0 @taps 0 0 16 112
// Retrieval info: CONNECT: taps80x 0 0 16 0 @taps 0 0 16 1280
// Retrieval info: CONNECT: taps81x 0 0 16 0 @taps 0 0 16 1296
// Retrieval info: CONNECT: taps82x 0 0 16 0 @taps 0 0 16 1312
// Retrieval info: CONNECT: taps83x 0 0 16 0 @taps 0 0 16 1328
// Retrieval info: CONNECT: taps84x 0 0 16 0 @taps 0 0 16 1344
// Retrieval info: CONNECT: taps85x 0 0 16 0 @taps 0 0 16 1360
// Retrieval info: CONNECT: taps86x 0 0 16 0 @taps 0 0 16 1376
// Retrieval info: CONNECT: taps87x 0 0 16 0 @taps 0 0 16 1392
// Retrieval info: CONNECT: taps88x 0 0 16 0 @taps 0 0 16 1408
// Retrieval info: CONNECT: taps89x 0 0 16 0 @taps 0 0 16 1424
// Retrieval info: CONNECT: taps8x 0 0 16 0 @taps 0 0 16 128
// Retrieval info: CONNECT: taps90x 0 0 16 0 @taps 0 0 16 1440
// Retrieval info: CONNECT: taps91x 0 0 16 0 @taps 0 0 16 1456
// Retrieval info: CONNECT: taps92x 0 0 16 0 @taps 0 0 16 1472
// Retrieval info: CONNECT: taps93x 0 0 16 0 @taps 0 0 16 1488
// Retrieval info: CONNECT: taps94x 0 0 16 0 @taps 0 0 16 1504
// Retrieval info: CONNECT: taps95x 0 0 16 0 @taps 0 0 16 1520
// Retrieval info: CONNECT: taps9x 0 0 16 0 @taps 0 0 16 144
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Shift_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
